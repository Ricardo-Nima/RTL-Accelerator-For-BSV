`timescale 1ns/1ns
module testbench();
 reg CLK, RST_N;
 reg [31 : 0] counter$count;
 reg  counter$overflow;
 mkTb U1(.CLK(CLK), 
		.RST_N(RST_N), 
		.counter$count(counter$count), 
		.counter$overflow(counter$overflow));
always begin
	#5 CLK = ~CLK;
end
initial begin
	RST_N = 0;
	#1 CLK = 1;
	#1 RST_N = 1;
end
 // port: counter$count
initial begin
	#0 counter$count = 18446744072277895850;
	#10 counter$count = 0;
	#10 counter$count = 1;
	#10 counter$count = 2;
	#10 counter$count = 3;
	#10 counter$count = 4;
	#10 counter$count = 5;
	#10 counter$count = 6;
	#10 counter$count = 7;
	#10 counter$count = 8;
	#10 counter$count = 9;
	#10 counter$count = 10;
	#10 counter$count = 11;
	#10 counter$count = 12;
	#10 counter$count = 13;
	#10 counter$count = 14;
	#10 counter$count = 15;
	#10 counter$count = 16;
	#10 counter$count = 17;
	#10 counter$count = 18;
	#10 counter$count = 19;
	#10 counter$count = 20;
	#10 counter$count = 21;
	#10 counter$count = 22;
	#10 counter$count = 23;
	#10 counter$count = 24;
	#10 counter$count = 25;
	#10 counter$count = 26;
	#10 counter$count = 27;
	#10 counter$count = 28;
	#10 counter$count = 29;
	#10 counter$count = 30;
	#10 counter$count = 31;
	#10 counter$count = 32;
	#10 counter$count = 33;
	#10 counter$count = 34;
	#10 counter$count = 35;
	#10 counter$count = 36;
	#10 counter$count = 37;
	#10 counter$count = 38;
	#10 counter$count = 39;
	#10 counter$count = 40;
	#10 counter$count = 41;
	#10 counter$count = 42;
	#10 counter$count = 43;
	#10 counter$count = 44;
	#10 counter$count = 45;
	#10 counter$count = 46;
	#10 counter$count = 47;
	#10 counter$count = 48;
	#10 counter$count = 49;
	#10 counter$count = 50;
	#10 counter$count = 51;
	#10 counter$count = 52;
	#10 counter$count = 53;
	#10 counter$count = 54;
	#10 counter$count = 55;
	#10 counter$count = 56;
	#10 counter$count = 57;
	#10 counter$count = 58;
	#10 counter$count = 59;
	#10 counter$count = 60;
	#10 counter$count = 61;
	#10 counter$count = 62;
	#10 counter$count = 63;
	#10 counter$count = 64;
	#10 counter$count = 65;
	#10 counter$count = 66;
	#10 counter$count = 67;
	#10 counter$count = 68;
	#10 counter$count = 69;
	#10 counter$count = 70;
	#10 counter$count = 71;
	#10 counter$count = 72;
	#10 counter$count = 73;
	#10 counter$count = 74;
	#10 counter$count = 75;
	#10 counter$count = 76;
	#10 counter$count = 77;
	#10 counter$count = 78;
	#10 counter$count = 79;
	#10 counter$count = 80;
	#10 counter$count = 81;
	#10 counter$count = 82;
	#10 counter$count = 83;
	#10 counter$count = 84;
	#10 counter$count = 85;
	#10 counter$count = 86;
	#10 counter$count = 87;
	#10 counter$count = 88;
	#10 counter$count = 89;
	#10 counter$count = 90;
	#10 counter$count = 91;
	#10 counter$count = 92;
	#10 counter$count = 93;
	#10 counter$count = 94;
	#10 counter$count = 95;
	#10 counter$count = 96;
	#10 counter$count = 97;
	#10 counter$count = 98;
	#10 counter$count = 99;
	#10 counter$count = 100;
	#10 counter$count = 101;
	#10 counter$count = 102;
	#10 counter$count = 103;
	#10 counter$count = 104;
	#10 counter$count = 105;
	#10 counter$count = 106;
	#10 counter$count = 107;
	#10 counter$count = 108;
	#10 counter$count = 109;
	#10 counter$count = 110;
	#10 counter$count = 111;
	#10 counter$count = 112;
	#10 counter$count = 113;
	#10 counter$count = 114;
	#10 counter$count = 115;
	#10 counter$count = 116;
	#10 counter$count = 117;
	#10 counter$count = 118;
	#10 counter$count = 119;
	#10 counter$count = 120;
	#10 counter$count = 121;
	#10 counter$count = 122;
	#10 counter$count = 123;
	#10 counter$count = 124;
	#10 counter$count = 125;
	#10 counter$count = 126;
	#10 counter$count = 127;
	#10 counter$count = 128;
	#10 counter$count = 129;
	#10 counter$count = 130;
	#10 counter$count = 131;
	#10 counter$count = 132;
	#10 counter$count = 133;
	#10 counter$count = 134;
	#10 counter$count = 135;
	#10 counter$count = 136;
	#10 counter$count = 137;
	#10 counter$count = 138;
	#10 counter$count = 139;
	#10 counter$count = 140;
	#10 counter$count = 141;
	#10 counter$count = 142;
	#10 counter$count = 143;
	#10 counter$count = 144;
	#10 counter$count = 145;
	#10 counter$count = 146;
	#10 counter$count = 147;
	#10 counter$count = 148;
	#10 counter$count = 149;
	#10 counter$count = 150;
	#10 counter$count = 151;
	#10 counter$count = 152;
	#10 counter$count = 153;
	#10 counter$count = 154;
	#10 counter$count = 155;
	#10 counter$count = 156;
	#10 counter$count = 157;
	#10 counter$count = 158;
	#10 counter$count = 159;
	#10 counter$count = 160;
	#10 counter$count = 161;
	#10 counter$count = 162;
	#10 counter$count = 163;
	#10 counter$count = 164;
	#10 counter$count = 165;
	#10 counter$count = 166;
	#10 counter$count = 167;
	#10 counter$count = 168;
	#10 counter$count = 169;
	#10 counter$count = 170;
	#10 counter$count = 171;
	#10 counter$count = 172;
	#10 counter$count = 173;
	#10 counter$count = 174;
	#10 counter$count = 175;
	#10 counter$count = 176;
	#10 counter$count = 177;
	#10 counter$count = 178;
	#10 counter$count = 179;
	#10 counter$count = 180;
	#10 counter$count = 181;
	#10 counter$count = 182;
	#10 counter$count = 183;
	#10 counter$count = 184;
	#10 counter$count = 185;
	#10 counter$count = 186;
	#10 counter$count = 187;
	#10 counter$count = 188;
	#10 counter$count = 189;
	#10 counter$count = 190;
	#10 counter$count = 191;
	#10 counter$count = 192;
	#10 counter$count = 193;
	#10 counter$count = 194;
	#10 counter$count = 195;
	#10 counter$count = 196;
	#10 counter$count = 197;
	#10 counter$count = 198;
	#10 counter$count = 199;
	#10 counter$count = 200;
	#10 counter$count = 201;
	#10 counter$count = 202;
	#10 counter$count = 203;
	#10 counter$count = 204;
	#10 counter$count = 205;
	#10 counter$count = 206;
	#10 counter$count = 207;
	#10 counter$count = 208;
	#10 counter$count = 209;
	#10 counter$count = 210;
	#10 counter$count = 211;
	#10 counter$count = 212;
	#10 counter$count = 213;
	#10 counter$count = 214;
	#10 counter$count = 215;
	#10 counter$count = 216;
	#10 counter$count = 217;
	#10 counter$count = 218;
	#10 counter$count = 219;
	#10 counter$count = 220;
	#10 counter$count = 221;
	#10 counter$count = 222;
	#10 counter$count = 223;
	#10 counter$count = 224;
	#10 counter$count = 225;
	#10 counter$count = 226;
	#10 counter$count = 227;
	#10 counter$count = 228;
	#10 counter$count = 229;
	#10 counter$count = 230;
	#10 counter$count = 231;
	#10 counter$count = 232;
	#10 counter$count = 233;
	#10 counter$count = 234;
	#10 counter$count = 235;
	#10 counter$count = 236;
	#10 counter$count = 237;
	#10 counter$count = 238;
	#10 counter$count = 239;
	#10 counter$count = 240;
	#10 counter$count = 241;
	#10 counter$count = 242;
	#10 counter$count = 243;
	#10 counter$count = 244;
	#10 counter$count = 245;
	#10 counter$count = 246;
	#10 counter$count = 247;
	#10 counter$count = 248;
	#10 counter$count = 249;
	#10 counter$count = 250;
	#10 counter$count = 251;
	#10 counter$count = 252;
	#10 counter$count = 253;
	#10 counter$count = 254;
	#10 counter$count = 255;
	#10 counter$count = 256;
	#10 counter$count = 257;
	#10 counter$count = 258;
	#10 counter$count = 259;
	#10 counter$count = 260;
	#10 counter$count = 261;
	#10 counter$count = 262;
	#10 counter$count = 263;
	#10 counter$count = 264;
	#10 counter$count = 265;
	#10 counter$count = 266;
	#10 counter$count = 267;
	#10 counter$count = 268;
	#10 counter$count = 269;
	#10 counter$count = 270;
	#10 counter$count = 271;
	#10 counter$count = 272;
	#10 counter$count = 273;
	#10 counter$count = 274;
	#10 counter$count = 275;
	#10 counter$count = 276;
	#10 counter$count = 277;
	#10 counter$count = 278;
	#10 counter$count = 279;
	#10 counter$count = 280;
	#10 counter$count = 281;
	#10 counter$count = 282;
	#10 counter$count = 283;
	#10 counter$count = 284;
	#10 counter$count = 285;
	#10 counter$count = 286;
	#10 counter$count = 287;
	#10 counter$count = 288;
	#10 counter$count = 289;
	#10 counter$count = 290;
	#10 counter$count = 291;
	#10 counter$count = 292;
	#10 counter$count = 293;
	#10 counter$count = 294;
	#10 counter$count = 295;
	#10 counter$count = 296;
	#10 counter$count = 297;
	#10 counter$count = 298;
	#10 counter$count = 299;
	#10 counter$count = 300;
	#10 counter$count = 301;
	#10 counter$count = 302;
	#10 counter$count = 303;
	#10 counter$count = 304;
	#10 counter$count = 305;
	#10 counter$count = 306;
	#10 counter$count = 307;
	#10 counter$count = 308;
	#10 counter$count = 309;
	#10 counter$count = 310;
	#10 counter$count = 311;
	#10 counter$count = 312;
	#10 counter$count = 313;
	#10 counter$count = 314;
	#10 counter$count = 315;
	#10 counter$count = 316;
	#10 counter$count = 317;
	#10 counter$count = 318;
	#10 counter$count = 319;
	#10 counter$count = 320;
	#10 counter$count = 321;
	#10 counter$count = 322;
	#10 counter$count = 323;
	#10 counter$count = 324;
	#10 counter$count = 325;
	#10 counter$count = 326;
	#10 counter$count = 327;
	#10 counter$count = 328;
	#10 counter$count = 329;
	#10 counter$count = 330;
	#10 counter$count = 331;
	#10 counter$count = 332;
	#10 counter$count = 333;
	#10 counter$count = 334;
	#10 counter$count = 335;
	#10 counter$count = 336;
	#10 counter$count = 337;
	#10 counter$count = 338;
	#10 counter$count = 339;
	#10 counter$count = 340;
	#10 counter$count = 341;
	#10 counter$count = 342;
	#10 counter$count = 343;
	#10 counter$count = 344;
	#10 counter$count = 345;
	#10 counter$count = 346;
	#10 counter$count = 347;
	#10 counter$count = 348;
	#10 counter$count = 349;
	#10 counter$count = 350;
	#10 counter$count = 351;
	#10 counter$count = 352;
	#10 counter$count = 353;
	#10 counter$count = 354;
	#10 counter$count = 355;
	#10 counter$count = 356;
	#10 counter$count = 357;
	#10 counter$count = 358;
	#10 counter$count = 359;
	#10 counter$count = 360;
	#10 counter$count = 361;
	#10 counter$count = 362;
	#10 counter$count = 363;
	#10 counter$count = 364;
	#10 counter$count = 365;
	#10 counter$count = 366;
	#10 counter$count = 367;
	#10 counter$count = 368;
	#10 counter$count = 369;
	#10 counter$count = 370;
	#10 counter$count = 371;
	#10 counter$count = 372;
	#10 counter$count = 373;
	#10 counter$count = 374;
	#10 counter$count = 375;
	#10 counter$count = 376;
	#10 counter$count = 377;
	#10 counter$count = 378;
	#10 counter$count = 379;
	#10 counter$count = 380;
	#10 counter$count = 381;
	#10 counter$count = 382;
	#10 counter$count = 383;
	#10 counter$count = 384;
	#10 counter$count = 385;
	#10 counter$count = 386;
	#10 counter$count = 387;
	#10 counter$count = 388;
	#10 counter$count = 389;
	#10 counter$count = 390;
	#10 counter$count = 391;
	#10 counter$count = 392;
	#10 counter$count = 393;
	#10 counter$count = 394;
	#10 counter$count = 395;
	#10 counter$count = 396;
	#10 counter$count = 397;
	#10 counter$count = 398;
	#10 counter$count = 399;
	#10 counter$count = 400;
	#10 counter$count = 401;
	#10 counter$count = 402;
	#10 counter$count = 403;
	#10 counter$count = 404;
	#10 counter$count = 405;
	#10 counter$count = 406;
	#10 counter$count = 407;
	#10 counter$count = 408;
	#10 counter$count = 409;
	#10 counter$count = 410;
	#10 counter$count = 411;
	#10 counter$count = 412;
	#10 counter$count = 413;
	#10 counter$count = 414;
	#10 counter$count = 415;
	#10 counter$count = 416;
	#10 counter$count = 417;
	#10 counter$count = 418;
	#10 counter$count = 419;
	#10 counter$count = 420;
	#10 counter$count = 421;
	#10 counter$count = 422;
	#10 counter$count = 423;
	#10 counter$count = 424;
	#10 counter$count = 425;
	#10 counter$count = 426;
	#10 counter$count = 427;
	#10 counter$count = 428;
	#10 counter$count = 429;
	#10 counter$count = 430;
	#10 counter$count = 431;
	#10 counter$count = 432;
	#10 counter$count = 433;
	#10 counter$count = 434;
	#10 counter$count = 435;
	#10 counter$count = 436;
	#10 counter$count = 437;
	#10 counter$count = 438;
	#10 counter$count = 439;
	#10 counter$count = 440;
	#10 counter$count = 441;
	#10 counter$count = 442;
	#10 counter$count = 443;
	#10 counter$count = 444;
	#10 counter$count = 445;
	#10 counter$count = 446;
	#10 counter$count = 447;
	#10 counter$count = 448;
	#10 counter$count = 449;
	#10 counter$count = 450;
	#10 counter$count = 451;
	#10 counter$count = 452;
	#10 counter$count = 453;
	#10 counter$count = 454;
	#10 counter$count = 455;
	#10 counter$count = 456;
	#10 counter$count = 457;
	#10 counter$count = 458;
	#10 counter$count = 459;
	#10 counter$count = 460;
	#10 counter$count = 461;
	#10 counter$count = 462;
	#10 counter$count = 463;
	#10 counter$count = 464;
	#10 counter$count = 465;
	#10 counter$count = 466;
	#10 counter$count = 467;
	#10 counter$count = 468;
	#10 counter$count = 469;
	#10 counter$count = 470;
	#10 counter$count = 471;
	#10 counter$count = 472;
	#10 counter$count = 473;
	#10 counter$count = 474;
	#10 counter$count = 475;
	#10 counter$count = 476;
	#10 counter$count = 477;
	#10 counter$count = 478;
	#10 counter$count = 479;
	#10 counter$count = 480;
	#10 counter$count = 481;
	#10 counter$count = 482;
	#10 counter$count = 483;
	#10 counter$count = 484;
	#10 counter$count = 485;
	#10 counter$count = 486;
	#10 counter$count = 487;
	#10 counter$count = 488;
	#10 counter$count = 489;
	#10 counter$count = 490;
	#10 counter$count = 491;
	#10 counter$count = 492;
	#10 counter$count = 493;
	#10 counter$count = 494;
	#10 counter$count = 495;
	#10 counter$count = 496;
	#10 counter$count = 497;
	#10 counter$count = 498;
	#10 counter$count = 499;
	#10 counter$count = 500;
	#10 counter$count = 501;
	#10 counter$count = 502;
	#10 counter$count = 503;
	#10 counter$count = 504;
	#10 counter$count = 505;
	#10 counter$count = 506;
	#10 counter$count = 507;
	#10 counter$count = 508;
	#10 counter$count = 509;
	#10 counter$count = 510;
	#10 counter$count = 511;
	#10 counter$count = 512;
	#10 counter$count = 513;
	#10 counter$count = 514;
	#10 counter$count = 515;
	#10 counter$count = 516;
	#10 counter$count = 517;
	#10 counter$count = 518;
	#10 counter$count = 519;
	#10 counter$count = 520;
	#10 counter$count = 521;
	#10 counter$count = 522;
	#10 counter$count = 523;
	#10 counter$count = 524;
	#10 counter$count = 525;
	#10 counter$count = 526;
	#10 counter$count = 527;
	#10 counter$count = 528;
	#10 counter$count = 529;
	#10 counter$count = 530;
	#10 counter$count = 531;
	#10 counter$count = 532;
	#10 counter$count = 533;
	#10 counter$count = 534;
	#10 counter$count = 535;
	#10 counter$count = 536;
	#10 counter$count = 537;
	#10 counter$count = 538;
	#10 counter$count = 539;
	#10 counter$count = 540;
	#10 counter$count = 541;
	#10 counter$count = 542;
	#10 counter$count = 543;
	#10 counter$count = 544;
	#10 counter$count = 545;
	#10 counter$count = 546;
	#10 counter$count = 547;
	#10 counter$count = 548;
	#10 counter$count = 549;
	#10 counter$count = 550;
	#10 counter$count = 551;
	#10 counter$count = 552;
	#10 counter$count = 553;
	#10 counter$count = 554;
	#10 counter$count = 555;
	#10 counter$count = 556;
	#10 counter$count = 557;
	#10 counter$count = 558;
	#10 counter$count = 559;
	#10 counter$count = 560;
	#10 counter$count = 561;
	#10 counter$count = 562;
	#10 counter$count = 563;
	#10 counter$count = 564;
	#10 counter$count = 565;
	#10 counter$count = 566;
	#10 counter$count = 567;
	#10 counter$count = 568;
	#10 counter$count = 569;
	#10 counter$count = 570;
	#10 counter$count = 571;
	#10 counter$count = 572;
	#10 counter$count = 573;
	#10 counter$count = 574;
	#10 counter$count = 575;
	#10 counter$count = 576;
	#10 counter$count = 577;
	#10 counter$count = 578;
	#10 counter$count = 579;
	#10 counter$count = 580;
	#10 counter$count = 581;
	#10 counter$count = 582;
	#10 counter$count = 583;
	#10 counter$count = 584;
	#10 counter$count = 585;
	#10 counter$count = 586;
	#10 counter$count = 587;
	#10 counter$count = 588;
	#10 counter$count = 589;
	#10 counter$count = 590;
	#10 counter$count = 591;
	#10 counter$count = 592;
	#10 counter$count = 593;
	#10 counter$count = 594;
	#10 counter$count = 595;
	#10 counter$count = 596;
	#10 counter$count = 597;
	#10 counter$count = 598;
	#10 counter$count = 599;
	#10 counter$count = 600;
	#10 counter$count = 601;
	#10 counter$count = 602;
	#10 counter$count = 603;
	#10 counter$count = 604;
	#10 counter$count = 605;
	#10 counter$count = 606;
	#10 counter$count = 607;
	#10 counter$count = 608;
	#10 counter$count = 609;
	#10 counter$count = 610;
	#10 counter$count = 611;
	#10 counter$count = 612;
	#10 counter$count = 613;
	#10 counter$count = 614;
	#10 counter$count = 615;
	#10 counter$count = 616;
	#10 counter$count = 617;
	#10 counter$count = 618;
	#10 counter$count = 619;
	#10 counter$count = 620;
	#10 counter$count = 621;
	#10 counter$count = 622;
	#10 counter$count = 623;
	#10 counter$count = 624;
	#10 counter$count = 625;
	#10 counter$count = 626;
	#10 counter$count = 627;
	#10 counter$count = 628;
	#10 counter$count = 629;
	#10 counter$count = 630;
	#10 counter$count = 631;
	#10 counter$count = 632;
	#10 counter$count = 633;
	#10 counter$count = 634;
	#10 counter$count = 635;
	#10 counter$count = 636;
	#10 counter$count = 637;
	#10 counter$count = 638;
	#10 counter$count = 639;
	#10 counter$count = 640;
	#10 counter$count = 641;
	#10 counter$count = 642;
	#10 counter$count = 643;
	#10 counter$count = 644;
	#10 counter$count = 645;
	#10 counter$count = 646;
	#10 counter$count = 647;
	#10 counter$count = 648;
	#10 counter$count = 649;
	#10 counter$count = 650;
	#10 counter$count = 651;
	#10 counter$count = 652;
	#10 counter$count = 653;
	#10 counter$count = 654;
	#10 counter$count = 655;
	#10 counter$count = 656;
	#10 counter$count = 657;
	#10 counter$count = 658;
	#10 counter$count = 659;
	#10 counter$count = 660;
	#10 counter$count = 661;
	#10 counter$count = 662;
	#10 counter$count = 663;
	#10 counter$count = 664;
	#10 counter$count = 665;
	#10 counter$count = 666;
	#10 counter$count = 667;
	#10 counter$count = 668;
	#10 counter$count = 669;
	#10 counter$count = 670;
	#10 counter$count = 671;
	#10 counter$count = 672;
	#10 counter$count = 673;
	#10 counter$count = 674;
	#10 counter$count = 675;
	#10 counter$count = 676;
	#10 counter$count = 677;
	#10 counter$count = 678;
	#10 counter$count = 679;
	#10 counter$count = 680;
	#10 counter$count = 681;
	#10 counter$count = 682;
	#10 counter$count = 683;
	#10 counter$count = 684;
	#10 counter$count = 685;
	#10 counter$count = 686;
	#10 counter$count = 687;
	#10 counter$count = 688;
	#10 counter$count = 689;
	#10 counter$count = 690;
	#10 counter$count = 691;
	#10 counter$count = 692;
	#10 counter$count = 693;
	#10 counter$count = 694;
	#10 counter$count = 695;
	#10 counter$count = 696;
	#10 counter$count = 697;
	#10 counter$count = 698;
	#10 counter$count = 699;
	#10 counter$count = 700;
	#10 counter$count = 701;
	#10 counter$count = 702;
	#10 counter$count = 703;
	#10 counter$count = 704;
	#10 counter$count = 705;
	#10 counter$count = 706;
	#10 counter$count = 707;
	#10 counter$count = 708;
	#10 counter$count = 709;
	#10 counter$count = 710;
	#10 counter$count = 711;
	#10 counter$count = 712;
	#10 counter$count = 713;
	#10 counter$count = 714;
	#10 counter$count = 715;
	#10 counter$count = 716;
	#10 counter$count = 717;
	#10 counter$count = 718;
	#10 counter$count = 719;
	#10 counter$count = 720;
	#10 counter$count = 721;
	#10 counter$count = 722;
	#10 counter$count = 723;
	#10 counter$count = 724;
	#10 counter$count = 725;
	#10 counter$count = 726;
	#10 counter$count = 727;
	#10 counter$count = 728;
	#10 counter$count = 729;
	#10 counter$count = 730;
	#10 counter$count = 731;
	#10 counter$count = 732;
	#10 counter$count = 733;
	#10 counter$count = 734;
	#10 counter$count = 735;
	#10 counter$count = 736;
	#10 counter$count = 737;
	#10 counter$count = 738;
	#10 counter$count = 739;
	#10 counter$count = 740;
	#10 counter$count = 741;
	#10 counter$count = 742;
	#10 counter$count = 743;
	#10 counter$count = 744;
	#10 counter$count = 745;
	#10 counter$count = 746;
	#10 counter$count = 747;
	#10 counter$count = 748;
	#10 counter$count = 749;
	#10 counter$count = 750;
	#10 counter$count = 751;
	#10 counter$count = 752;
	#10 counter$count = 753;
	#10 counter$count = 754;
	#10 counter$count = 755;
	#10 counter$count = 756;
	#10 counter$count = 757;
	#10 counter$count = 758;
	#10 counter$count = 759;
	#10 counter$count = 760;
	#10 counter$count = 761;
	#10 counter$count = 762;
	#10 counter$count = 763;
	#10 counter$count = 764;
	#10 counter$count = 765;
	#10 counter$count = 766;
	#10 counter$count = 767;
	#10 counter$count = 768;
	#10 counter$count = 769;
	#10 counter$count = 770;
	#10 counter$count = 771;
	#10 counter$count = 772;
	#10 counter$count = 773;
	#10 counter$count = 774;
	#10 counter$count = 775;
	#10 counter$count = 776;
	#10 counter$count = 777;
	#10 counter$count = 778;
	#10 counter$count = 779;
	#10 counter$count = 780;
	#10 counter$count = 781;
	#10 counter$count = 782;
	#10 counter$count = 783;
	#10 counter$count = 784;
	#10 counter$count = 785;
	#10 counter$count = 786;
	#10 counter$count = 787;
	#10 counter$count = 788;
	#10 counter$count = 789;
	#10 counter$count = 790;
	#10 counter$count = 791;
	#10 counter$count = 792;
	#10 counter$count = 793;
	#10 counter$count = 794;
	#10 counter$count = 795;
	#10 counter$count = 796;
	#10 counter$count = 797;
	#10 counter$count = 798;
	#10 counter$count = 799;
	#10 counter$count = 800;
	#10 counter$count = 801;
	#10 counter$count = 802;
	#10 counter$count = 803;
	#10 counter$count = 804;
	#10 counter$count = 805;
	#10 counter$count = 806;
	#10 counter$count = 807;
	#10 counter$count = 808;
	#10 counter$count = 809;
	#10 counter$count = 810;
	#10 counter$count = 811;
	#10 counter$count = 812;
	#10 counter$count = 813;
	#10 counter$count = 814;
	#10 counter$count = 815;
	#10 counter$count = 816;
	#10 counter$count = 817;
	#10 counter$count = 818;
	#10 counter$count = 819;
	#10 counter$count = 820;
	#10 counter$count = 821;
	#10 counter$count = 822;
	#10 counter$count = 823;
	#10 counter$count = 824;
	#10 counter$count = 825;
	#10 counter$count = 826;
	#10 counter$count = 827;
	#10 counter$count = 828;
	#10 counter$count = 829;
	#10 counter$count = 830;
	#10 counter$count = 831;
	#10 counter$count = 832;
	#10 counter$count = 833;
	#10 counter$count = 834;
	#10 counter$count = 835;
	#10 counter$count = 836;
	#10 counter$count = 837;
	#10 counter$count = 838;
	#10 counter$count = 839;
	#10 counter$count = 840;
	#10 counter$count = 841;
	#10 counter$count = 842;
	#10 counter$count = 843;
	#10 counter$count = 844;
	#10 counter$count = 845;
	#10 counter$count = 846;
	#10 counter$count = 847;
	#10 counter$count = 848;
	#10 counter$count = 849;
	#10 counter$count = 850;
	#10 counter$count = 851;
	#10 counter$count = 852;
	#10 counter$count = 853;
	#10 counter$count = 854;
	#10 counter$count = 855;
	#10 counter$count = 856;
	#10 counter$count = 857;
	#10 counter$count = 858;
	#10 counter$count = 859;
	#10 counter$count = 860;
	#10 counter$count = 861;
	#10 counter$count = 862;
	#10 counter$count = 863;
	#10 counter$count = 864;
	#10 counter$count = 865;
	#10 counter$count = 866;
	#10 counter$count = 867;
	#10 counter$count = 868;
	#10 counter$count = 869;
	#10 counter$count = 870;
	#10 counter$count = 871;
	#10 counter$count = 872;
	#10 counter$count = 873;
	#10 counter$count = 874;
	#10 counter$count = 875;
	#10 counter$count = 876;
	#10 counter$count = 877;
	#10 counter$count = 878;
	#10 counter$count = 879;
	#10 counter$count = 880;
	#10 counter$count = 881;
	#10 counter$count = 882;
	#10 counter$count = 883;
	#10 counter$count = 884;
	#10 counter$count = 885;
	#10 counter$count = 886;
	#10 counter$count = 887;
	#10 counter$count = 888;
	#10 counter$count = 889;
	#10 counter$count = 890;
	#10 counter$count = 891;
	#10 counter$count = 892;
	#10 counter$count = 893;
	#10 counter$count = 894;
	#10 counter$count = 895;
	#10 counter$count = 896;
	#10 counter$count = 897;
	#10 counter$count = 898;
	#10 counter$count = 899;
	#10 counter$count = 900;
	#10 counter$count = 901;
	#10 counter$count = 902;
	#10 counter$count = 903;
	#10 counter$count = 904;
	#10 counter$count = 905;
	#10 counter$count = 906;
	#10 counter$count = 907;
	#10 counter$count = 908;
	#10 counter$count = 909;
	#10 counter$count = 910;
	#10 counter$count = 911;
	#10 counter$count = 912;
	#10 counter$count = 913;
	#10 counter$count = 914;
	#10 counter$count = 915;
	#10 counter$count = 916;
	#10 counter$count = 917;
	#10 counter$count = 918;
	#10 counter$count = 919;
	#10 counter$count = 920;
	#10 counter$count = 921;
	#10 counter$count = 922;
	#10 counter$count = 923;
	#10 counter$count = 924;
	#10 counter$count = 925;
	#10 counter$count = 926;
	#10 counter$count = 927;
	#10 counter$count = 928;
	#10 counter$count = 929;
	#10 counter$count = 930;
	#10 counter$count = 931;
	#10 counter$count = 932;
	#10 counter$count = 933;
	#10 counter$count = 934;
	#10 counter$count = 935;
	#10 counter$count = 936;
	#10 counter$count = 937;
	#10 counter$count = 938;
	#10 counter$count = 939;
	#10 counter$count = 940;
	#10 counter$count = 941;
	#10 counter$count = 942;
	#10 counter$count = 943;
	#10 counter$count = 944;
	#10 counter$count = 945;
	#10 counter$count = 946;
	#10 counter$count = 947;
	#10 counter$count = 948;
	#10 counter$count = 949;
	#10 counter$count = 950;
	#10 counter$count = 951;
	#10 counter$count = 952;
	#10 counter$count = 953;
	#10 counter$count = 954;
	#10 counter$count = 955;
	#10 counter$count = 956;
	#10 counter$count = 957;
	#10 counter$count = 958;
	#10 counter$count = 959;
	#10 counter$count = 960;
	#10 counter$count = 961;
	#10 counter$count = 962;
	#10 counter$count = 963;
	#10 counter$count = 964;
	#10 counter$count = 965;
	#10 counter$count = 966;
	#10 counter$count = 967;
	#10 counter$count = 968;
	#10 counter$count = 969;
	#10 counter$count = 970;
	#10 counter$count = 971;
	#10 counter$count = 972;
	#10 counter$count = 973;
	#10 counter$count = 974;
	#10 counter$count = 975;
	#10 counter$count = 976;
	#10 counter$count = 977;
	#10 counter$count = 978;
	#10 counter$count = 979;
	#10 counter$count = 980;
	#10 counter$count = 981;
	#10 counter$count = 982;
	#10 counter$count = 983;
	#10 counter$count = 984;
	#10 counter$count = 985;
	#10 counter$count = 986;
	#10 counter$count = 987;
	#10 counter$count = 988;
	#10 counter$count = 989;
	#10 counter$count = 990;
	#10 counter$count = 991;
	#10 counter$count = 992;
	#10 counter$count = 993;
	#10 counter$count = 994;
	#10 counter$count = 995;
	#10 counter$count = 996;
	#10 counter$count = 997;
	#10 counter$count = 998;
	#10 counter$count = 999;
	#10 counter$count = 1000;
	#10 counter$count = 1001;
	#10 counter$count = 1002;
	#10 counter$count = 1003;
	#10 counter$count = 1004;
	#10 counter$count = 1005;
	#10 counter$count = 1006;
	#10 counter$count = 1007;
	#10 counter$count = 1008;
	#10 counter$count = 1009;
	#10 counter$count = 1010;
	#10 counter$count = 1011;
	#10 counter$count = 1012;
	#10 counter$count = 1013;
	#10 counter$count = 1014;
	#10 counter$count = 1015;
	#10 counter$count = 1016;
	#10 counter$count = 1017;
	#10 counter$count = 1018;
	#10 counter$count = 1019;
	#10 counter$count = 1020;
	#10 counter$count = 1021;
	#10 counter$count = 1022;
	#10 counter$count = 1023;
	#10 counter$count = 1024;
	#10 counter$count = 1025;
	#10 counter$count = 1026;
	#10 counter$count = 1027;
	#10 counter$count = 1028;
	#10 counter$count = 1029;
	#10 counter$count = 1030;
	#10 counter$count = 1031;
	#10 counter$count = 1032;
	#10 counter$count = 1033;
	#10 counter$count = 1034;
	#10 counter$count = 1035;
	#10 counter$count = 1036;
	#10 counter$count = 1037;
	#10 counter$count = 1038;
	#10 counter$count = 1039;
	#10 counter$count = 1040;
	#10 counter$count = 1041;
	#10 counter$count = 1042;
	#10 counter$count = 1043;
	#10 counter$count = 1044;
	#10 counter$count = 1045;
	#10 counter$count = 1046;
	#10 counter$count = 1047;
	#10 counter$count = 1048;
	#10 counter$count = 1049;
	#10 counter$count = 1050;
	#10 counter$count = 1051;
	#10 counter$count = 1052;
	#10 counter$count = 1053;
	#10 counter$count = 1054;
	#10 counter$count = 1055;
	#10 counter$count = 1056;
	#10 counter$count = 1057;
	#10 counter$count = 1058;
	#10 counter$count = 1059;
	#10 counter$count = 1060;
	#10 counter$count = 1061;
	#10 counter$count = 1062;
	#10 counter$count = 1063;
	#10 counter$count = 1064;
	#10 counter$count = 1065;
	#10 counter$count = 1066;
	#10 counter$count = 1067;
	#10 counter$count = 1068;
	#10 counter$count = 1069;
	#10 counter$count = 1070;
	#10 counter$count = 1071;
	#10 counter$count = 1072;
	#10 counter$count = 1073;
	#10 counter$count = 1074;
	#10 counter$count = 1075;
	#10 counter$count = 1076;
	#10 counter$count = 1077;
	#10 counter$count = 1078;
	#10 counter$count = 1079;
	#10 counter$count = 1080;
	#10 counter$count = 1081;
	#10 counter$count = 1082;
	#10 counter$count = 1083;
	#10 counter$count = 1084;
	#10 counter$count = 1085;
	#10 counter$count = 1086;
	#10 counter$count = 1087;
	#10 counter$count = 1088;
	#10 counter$count = 1089;
	#10 counter$count = 1090;
	#10 counter$count = 1091;
	#10 counter$count = 1092;
	#10 counter$count = 1093;
	#10 counter$count = 1094;
	#10 counter$count = 1095;
	#10 counter$count = 1096;
	#10 counter$count = 1097;
	#10 counter$count = 1098;
	#10 counter$count = 1099;
	#10 counter$count = 1100;
	#10 counter$count = 1101;
	#10 counter$count = 1102;
	#10 counter$count = 1103;
	#10 counter$count = 1104;
	#10 counter$count = 1105;
	#10 counter$count = 1106;
	#10 counter$count = 1107;
	#10 counter$count = 1108;
	#10 counter$count = 1109;
	#10 counter$count = 1110;
	#10 counter$count = 1111;
	#10 counter$count = 1112;
	#10 counter$count = 1113;
	#10 counter$count = 1114;
	#10 counter$count = 1115;
	#10 counter$count = 1116;
	#10 counter$count = 1117;
	#10 counter$count = 1118;
	#10 counter$count = 1119;
	#10 counter$count = 1120;
	#10 counter$count = 1121;
	#10 counter$count = 1122;
	#10 counter$count = 1123;
	#10 counter$count = 1124;
	#10 counter$count = 1125;
	#10 counter$count = 1126;
	#10 counter$count = 1127;
	#10 counter$count = 1128;
	#10 counter$count = 1129;
	#10 counter$count = 1130;
	#10 counter$count = 1131;
	#10 counter$count = 1132;
	#10 counter$count = 1133;
	#10 counter$count = 1134;
	#10 counter$count = 1135;
	#10 counter$count = 1136;
	#10 counter$count = 1137;
	#10 counter$count = 1138;
	#10 counter$count = 1139;
	#10 counter$count = 1140;
	#10 counter$count = 1141;
	#10 counter$count = 1142;
	#10 counter$count = 1143;
	#10 counter$count = 1144;
	#10 counter$count = 1145;
	#10 counter$count = 1146;
	#10 counter$count = 1147;
	#10 counter$count = 1148;
	#10 counter$count = 1149;
	#10 counter$count = 1150;
	#10 counter$count = 1151;
	#10 counter$count = 1152;
	#10 counter$count = 1153;
	#10 counter$count = 1154;
	#10 counter$count = 1155;
	#10 counter$count = 1156;
	#10 counter$count = 1157;
	#10 counter$count = 1158;
	#10 counter$count = 1159;
	#10 counter$count = 1160;
	#10 counter$count = 1161;
	#10 counter$count = 1162;
	#10 counter$count = 1163;
	#10 counter$count = 1164;
	#10 counter$count = 1165;
	#10 counter$count = 1166;
	#10 counter$count = 1167;
	#10 counter$count = 1168;
	#10 counter$count = 1169;
	#10 counter$count = 1170;
	#10 counter$count = 1171;
	#10 counter$count = 1172;
	#10 counter$count = 1173;
	#10 counter$count = 1174;
	#10 counter$count = 1175;
	#10 counter$count = 1176;
	#10 counter$count = 1177;
	#10 counter$count = 1178;
	#10 counter$count = 1179;
	#10 counter$count = 1180;
	#10 counter$count = 1181;
	#10 counter$count = 1182;
	#10 counter$count = 1183;
	#10 counter$count = 1184;
	#10 counter$count = 1185;
	#10 counter$count = 1186;
	#10 counter$count = 1187;
	#10 counter$count = 1188;
	#10 counter$count = 1189;
	#10 counter$count = 1190;
	#10 counter$count = 1191;
	#10 counter$count = 1192;
	#10 counter$count = 1193;
	#10 counter$count = 1194;
	#10 counter$count = 1195;
	#10 counter$count = 1196;
	#10 counter$count = 1197;
	#10 counter$count = 1198;
	#10 counter$count = 1199;
	#10 counter$count = 1200;
	#10 counter$count = 1201;
	#10 counter$count = 1202;
	#10 counter$count = 1203;
	#10 counter$count = 1204;
	#10 counter$count = 1205;
	#10 counter$count = 1206;
	#10 counter$count = 1207;
	#10 counter$count = 1208;
	#10 counter$count = 1209;
	#10 counter$count = 1210;
	#10 counter$count = 1211;
	#10 counter$count = 1212;
	#10 counter$count = 1213;
	#10 counter$count = 1214;
	#10 counter$count = 1215;
	#10 counter$count = 1216;
	#10 counter$count = 1217;
	#10 counter$count = 1218;
	#10 counter$count = 1219;
	#10 counter$count = 1220;
	#10 counter$count = 1221;
	#10 counter$count = 1222;
	#10 counter$count = 1223;
	#10 counter$count = 1224;
	#10 counter$count = 1225;
	#10 counter$count = 1226;
	#10 counter$count = 1227;
	#10 counter$count = 1228;
	#10 counter$count = 1229;
	#10 counter$count = 1230;
	#10 counter$count = 1231;
	#10 counter$count = 1232;
	#10 counter$count = 1233;
	#10 counter$count = 1234;
	#10 counter$count = 1235;
	#10 counter$count = 1236;
	#10 counter$count = 1237;
	#10 counter$count = 1238;
	#10 counter$count = 1239;
	#10 counter$count = 1240;
	#10 counter$count = 1241;
	#10 counter$count = 1242;
	#10 counter$count = 1243;
	#10 counter$count = 1244;
	#10 counter$count = 1245;
	#10 counter$count = 1246;
	#10 counter$count = 1247;
	#10 counter$count = 1248;
	#10 counter$count = 1249;
	#10 counter$count = 1250;
	#10 counter$count = 1251;
	#10 counter$count = 1252;
	#10 counter$count = 1253;
	#10 counter$count = 1254;
	#10 counter$count = 1255;
	#10 counter$count = 1256;
	#10 counter$count = 1257;
	#10 counter$count = 1258;
	#10 counter$count = 1259;
	#10 counter$count = 1260;
	#10 counter$count = 1261;
	#10 counter$count = 1262;
	#10 counter$count = 1263;
	#10 counter$count = 1264;
	#10 counter$count = 1265;
	#10 counter$count = 1266;
	#10 counter$count = 1267;
	#10 counter$count = 1268;
	#10 counter$count = 1269;
	#10 counter$count = 1270;
	#10 counter$count = 1271;
	#10 counter$count = 1272;
	#10 counter$count = 1273;
	#10 counter$count = 1274;
	#10 counter$count = 1275;
	#10 counter$count = 1276;
	#10 counter$count = 1277;
	#10 counter$count = 1278;
	#10 counter$count = 1279;
	#10 counter$count = 1280;
	#10 counter$count = 1281;
	#10 counter$count = 1282;
	#10 counter$count = 1283;
	#10 counter$count = 1284;
	#10 counter$count = 1285;
	#10 counter$count = 1286;
	#10 counter$count = 1287;
	#10 counter$count = 1288;
	#10 counter$count = 1289;
	#10 counter$count = 1290;
	#10 counter$count = 1291;
	#10 counter$count = 1292;
	#10 counter$count = 1293;
	#10 counter$count = 1294;
	#10 counter$count = 1295;
	#10 counter$count = 1296;
	#10 counter$count = 1297;
	#10 counter$count = 1298;
	#10 counter$count = 1299;
	#10 counter$count = 1300;
	#10 counter$count = 1301;
	#10 counter$count = 1302;
	#10 counter$count = 1303;
	#10 counter$count = 1304;
	#10 counter$count = 1305;
	#10 counter$count = 1306;
	#10 counter$count = 1307;
	#10 counter$count = 1308;
	#10 counter$count = 1309;
	#10 counter$count = 1310;
	#10 counter$count = 1311;
	#10 counter$count = 1312;
	#10 counter$count = 1313;
	#10 counter$count = 1314;
	#10 counter$count = 1315;
	#10 counter$count = 1316;
	#10 counter$count = 1317;
	#10 counter$count = 1318;
	#10 counter$count = 1319;
	#10 counter$count = 1320;
	#10 counter$count = 1321;
	#10 counter$count = 1322;
	#10 counter$count = 1323;
	#10 counter$count = 1324;
	#10 counter$count = 1325;
	#10 counter$count = 1326;
	#10 counter$count = 1327;
	#10 counter$count = 1328;
	#10 counter$count = 1329;
	#10 counter$count = 1330;
	#10 counter$count = 1331;
	#10 counter$count = 1332;
	#10 counter$count = 1333;
	#10 counter$count = 1334;
	#10 counter$count = 1335;
	#10 counter$count = 1336;
	#10 counter$count = 1337;
	#10 counter$count = 1338;
	#10 counter$count = 1339;
	#10 counter$count = 1340;
	#10 counter$count = 1341;
	#10 counter$count = 1342;
	#10 counter$count = 1343;
	#10 counter$count = 1344;
	#10 counter$count = 1345;
	#10 counter$count = 1346;
	#10 counter$count = 1347;
	#10 counter$count = 1348;
	#10 counter$count = 1349;
	#10 counter$count = 1350;
	#10 counter$count = 1351;
	#10 counter$count = 1352;
	#10 counter$count = 1353;
	#10 counter$count = 1354;
	#10 counter$count = 1355;
	#10 counter$count = 1356;
	#10 counter$count = 1357;
	#10 counter$count = 1358;
	#10 counter$count = 1359;
	#10 counter$count = 1360;
	#10 counter$count = 1361;
	#10 counter$count = 1362;
	#10 counter$count = 1363;
	#10 counter$count = 1364;
	#10 counter$count = 1365;
	#10 counter$count = 1366;
	#10 counter$count = 1367;
	#10 counter$count = 1368;
	#10 counter$count = 1369;
	#10 counter$count = 1370;
	#10 counter$count = 1371;
	#10 counter$count = 1372;
	#10 counter$count = 1373;
	#10 counter$count = 1374;
	#10 counter$count = 1375;
	#10 counter$count = 1376;
	#10 counter$count = 1377;
	#10 counter$count = 1378;
	#10 counter$count = 1379;
	#10 counter$count = 1380;
	#10 counter$count = 1381;
	#10 counter$count = 1382;
	#10 counter$count = 1383;
	#10 counter$count = 1384;
	#10 counter$count = 1385;
	#10 counter$count = 1386;
	#10 counter$count = 1387;
	#10 counter$count = 1388;
	#10 counter$count = 1389;
	#10 counter$count = 1390;
	#10 counter$count = 1391;
	#10 counter$count = 1392;
	#10 counter$count = 1393;
	#10 counter$count = 1394;
	#10 counter$count = 1395;
	#10 counter$count = 1396;
	#10 counter$count = 1397;
	#10 counter$count = 1398;
	#10 counter$count = 1399;
	#10 counter$count = 1400;
	#10 counter$count = 1401;
	#10 counter$count = 1402;
	#10 counter$count = 1403;
	#10 counter$count = 1404;
	#10 counter$count = 1405;
	#10 counter$count = 1406;
	#10 counter$count = 1407;
	#10 counter$count = 1408;
	#10 counter$count = 1409;
	#10 counter$count = 1410;
	#10 counter$count = 1411;
	#10 counter$count = 1412;
	#10 counter$count = 1413;
	#10 counter$count = 1414;
	#10 counter$count = 1415;
	#10 counter$count = 1416;
	#10 counter$count = 1417;
	#10 counter$count = 1418;
	#10 counter$count = 1419;
	#10 counter$count = 1420;
	#10 counter$count = 1421;
	#10 counter$count = 1422;
	#10 counter$count = 1423;
	#10 counter$count = 1424;
	#10 counter$count = 1425;
	#10 counter$count = 1426;
	#10 counter$count = 1427;
	#10 counter$count = 1428;
	#10 counter$count = 1429;
	#10 counter$count = 1430;
	#10 counter$count = 1431;
	#10 counter$count = 1432;
	#10 counter$count = 1433;
	#10 counter$count = 1434;
	#10 counter$count = 1435;
	#10 counter$count = 1436;
	#10 counter$count = 1437;
	#10 counter$count = 1438;
	#10 counter$count = 1439;
	#10 counter$count = 1440;
	#10 counter$count = 1441;
	#10 counter$count = 1442;
	#10 counter$count = 1443;
	#10 counter$count = 1444;
	#10 counter$count = 1445;
	#10 counter$count = 1446;
	#10 counter$count = 1447;
	#10 counter$count = 1448;
	#10 counter$count = 1449;
	#10 counter$count = 1450;
	#10 counter$count = 1451;
	#10 counter$count = 1452;
	#10 counter$count = 1453;
	#10 counter$count = 1454;
	#10 counter$count = 1455;
	#10 counter$count = 1456;
	#10 counter$count = 1457;
	#10 counter$count = 1458;
	#10 counter$count = 1459;
	#10 counter$count = 1460;
	#10 counter$count = 1461;
	#10 counter$count = 1462;
	#10 counter$count = 1463;
	#10 counter$count = 1464;
	#10 counter$count = 1465;
	#10 counter$count = 1466;
	#10 counter$count = 1467;
	#10 counter$count = 1468;
	#10 counter$count = 1469;
	#10 counter$count = 1470;
	#10 counter$count = 1471;
	#10 counter$count = 1472;
	#10 counter$count = 1473;
	#10 counter$count = 1474;
	#10 counter$count = 1475;
	#10 counter$count = 1476;
	#10 counter$count = 1477;
	#10 counter$count = 1478;
	#10 counter$count = 1479;
	#10 counter$count = 1480;
	#10 counter$count = 1481;
	#10 counter$count = 1482;
	#10 counter$count = 1483;
	#10 counter$count = 1484;
	#10 counter$count = 1485;
	#10 counter$count = 1486;
	#10 counter$count = 1487;
	#10 counter$count = 1488;
	#10 counter$count = 1489;
	#10 counter$count = 1490;
	#10 counter$count = 1491;
	#10 counter$count = 1492;
	#10 counter$count = 1493;
	#10 counter$count = 1494;
	#10 counter$count = 1495;
	#10 counter$count = 1496;
	#10 counter$count = 1497;
	#10 counter$count = 1498;
	#10 counter$count = 1499;
	#10 counter$count = 1500;
	#10 counter$count = 1501;
	#10 counter$count = 1502;
	#10 counter$count = 1503;
	#10 counter$count = 1504;
	#10 counter$count = 1505;
	#10 counter$count = 1506;
	#10 counter$count = 1507;
	#10 counter$count = 1508;
	#10 counter$count = 1509;
	#10 counter$count = 1510;
	#10 counter$count = 1511;
	#10 counter$count = 1512;
	#10 counter$count = 1513;
	#10 counter$count = 1514;
	#10 counter$count = 1515;
	#10 counter$count = 1516;
	#10 counter$count = 1517;
	#10 counter$count = 1518;
	#10 counter$count = 1519;
	#10 counter$count = 1520;
	#10 counter$count = 1521;
	#10 counter$count = 1522;
	#10 counter$count = 1523;
	#10 counter$count = 1524;
	#10 counter$count = 1525;
	#10 counter$count = 1526;
	#10 counter$count = 1527;
	#10 counter$count = 1528;
	#10 counter$count = 1529;
	#10 counter$count = 1530;
	#10 counter$count = 1531;
	#10 counter$count = 1532;
	#10 counter$count = 1533;
	#10 counter$count = 1534;
	#10 counter$count = 1535;
	#10 counter$count = 1536;
	#10 counter$count = 1537;
	#10 counter$count = 1538;
	#10 counter$count = 1539;
	#10 counter$count = 1540;
	#10 counter$count = 1541;
	#10 counter$count = 1542;
	#10 counter$count = 1543;
	#10 counter$count = 1544;
	#10 counter$count = 1545;
	#10 counter$count = 1546;
	#10 counter$count = 1547;
	#10 counter$count = 1548;
	#10 counter$count = 1549;
	#10 counter$count = 1550;
	#10 counter$count = 1551;
	#10 counter$count = 1552;
	#10 counter$count = 1553;
	#10 counter$count = 1554;
	#10 counter$count = 1555;
	#10 counter$count = 1556;
	#10 counter$count = 1557;
	#10 counter$count = 1558;
	#10 counter$count = 1559;
	#10 counter$count = 1560;
	#10 counter$count = 1561;
	#10 counter$count = 1562;
	#10 counter$count = 1563;
	#10 counter$count = 1564;
	#10 counter$count = 1565;
	#10 counter$count = 1566;
	#10 counter$count = 1567;
	#10 counter$count = 1568;
	#10 counter$count = 1569;
	#10 counter$count = 1570;
	#10 counter$count = 1571;
	#10 counter$count = 1572;
	#10 counter$count = 1573;
	#10 counter$count = 1574;
	#10 counter$count = 1575;
	#10 counter$count = 1576;
	#10 counter$count = 1577;
	#10 counter$count = 1578;
	#10 counter$count = 1579;
	#10 counter$count = 1580;
	#10 counter$count = 1581;
	#10 counter$count = 1582;
	#10 counter$count = 1583;
	#10 counter$count = 1584;
	#10 counter$count = 1585;
	#10 counter$count = 1586;
	#10 counter$count = 1587;
	#10 counter$count = 1588;
	#10 counter$count = 1589;
	#10 counter$count = 1590;
	#10 counter$count = 1591;
	#10 counter$count = 1592;
	#10 counter$count = 1593;
	#10 counter$count = 1594;
	#10 counter$count = 1595;
	#10 counter$count = 1596;
	#10 counter$count = 1597;
	#10 counter$count = 1598;
	#10 counter$count = 1599;
	#10 counter$count = 1600;
	#10 counter$count = 1601;
	#10 counter$count = 1602;
	#10 counter$count = 1603;
	#10 counter$count = 1604;
	#10 counter$count = 1605;
	#10 counter$count = 1606;
	#10 counter$count = 1607;
	#10 counter$count = 1608;
	#10 counter$count = 1609;
	#10 counter$count = 1610;
	#10 counter$count = 1611;
	#10 counter$count = 1612;
	#10 counter$count = 1613;
	#10 counter$count = 1614;
	#10 counter$count = 1615;
	#10 counter$count = 1616;
	#10 counter$count = 1617;
	#10 counter$count = 1618;
	#10 counter$count = 1619;
	#10 counter$count = 1620;
	#10 counter$count = 1621;
	#10 counter$count = 1622;
	#10 counter$count = 1623;
	#10 counter$count = 1624;
	#10 counter$count = 1625;
	#10 counter$count = 1626;
	#10 counter$count = 1627;
	#10 counter$count = 1628;
	#10 counter$count = 1629;
	#10 counter$count = 1630;
	#10 counter$count = 1631;
	#10 counter$count = 1632;
	#10 counter$count = 1633;
	#10 counter$count = 1634;
	#10 counter$count = 1635;
	#10 counter$count = 1636;
	#10 counter$count = 1637;
	#10 counter$count = 1638;
	#10 counter$count = 1639;
	#10 counter$count = 1640;
	#10 counter$count = 1641;
	#10 counter$count = 1642;
	#10 counter$count = 1643;
	#10 counter$count = 1644;
	#10 counter$count = 1645;
	#10 counter$count = 1646;
	#10 counter$count = 1647;
	#10 counter$count = 1648;
	#10 counter$count = 1649;
	#10 counter$count = 1650;
	#10 counter$count = 1651;
	#10 counter$count = 1652;
	#10 counter$count = 1653;
	#10 counter$count = 1654;
	#10 counter$count = 1655;
	#10 counter$count = 1656;
	#10 counter$count = 1657;
	#10 counter$count = 1658;
	#10 counter$count = 1659;
	#10 counter$count = 1660;
	#10 counter$count = 1661;
	#10 counter$count = 1662;
	#10 counter$count = 1663;
	#10 counter$count = 1664;
	#10 counter$count = 1665;
	#10 counter$count = 1666;
	#10 counter$count = 1667;
	#10 counter$count = 1668;
	#10 counter$count = 1669;
	#10 counter$count = 1670;
	#10 counter$count = 1671;
	#10 counter$count = 1672;
	#10 counter$count = 1673;
	#10 counter$count = 1674;
	#10 counter$count = 1675;
	#10 counter$count = 1676;
	#10 counter$count = 1677;
	#10 counter$count = 1678;
	#10 counter$count = 1679;
	#10 counter$count = 1680;
	#10 counter$count = 1681;
	#10 counter$count = 1682;
	#10 counter$count = 1683;
	#10 counter$count = 1684;
	#10 counter$count = 1685;
	#10 counter$count = 1686;
	#10 counter$count = 1687;
	#10 counter$count = 1688;
	#10 counter$count = 1689;
	#10 counter$count = 1690;
	#10 counter$count = 1691;
	#10 counter$count = 1692;
	#10 counter$count = 1693;
	#10 counter$count = 1694;
	#10 counter$count = 1695;
	#10 counter$count = 1696;
	#10 counter$count = 1697;
	#10 counter$count = 1698;
	#10 counter$count = 1699;
	#10 counter$count = 1700;
	#10 counter$count = 1701;
	#10 counter$count = 1702;
	#10 counter$count = 1703;
	#10 counter$count = 1704;
	#10 counter$count = 1705;
	#10 counter$count = 1706;
	#10 counter$count = 1707;
	#10 counter$count = 1708;
	#10 counter$count = 1709;
	#10 counter$count = 1710;
	#10 counter$count = 1711;
	#10 counter$count = 1712;
	#10 counter$count = 1713;
	#10 counter$count = 1714;
	#10 counter$count = 1715;
	#10 counter$count = 1716;
	#10 counter$count = 1717;
	#10 counter$count = 1718;
	#10 counter$count = 1719;
	#10 counter$count = 1720;
	#10 counter$count = 1721;
	#10 counter$count = 1722;
	#10 counter$count = 1723;
	#10 counter$count = 1724;
	#10 counter$count = 1725;
	#10 counter$count = 1726;
	#10 counter$count = 1727;
	#10 counter$count = 1728;
	#10 counter$count = 1729;
	#10 counter$count = 1730;
	#10 counter$count = 1731;
	#10 counter$count = 1732;
	#10 counter$count = 1733;
	#10 counter$count = 1734;
	#10 counter$count = 1735;
	#10 counter$count = 1736;
	#10 counter$count = 1737;
	#10 counter$count = 1738;
	#10 counter$count = 1739;
	#10 counter$count = 1740;
	#10 counter$count = 1741;
	#10 counter$count = 1742;
	#10 counter$count = 1743;
	#10 counter$count = 1744;
	#10 counter$count = 1745;
	#10 counter$count = 1746;
	#10 counter$count = 1747;
	#10 counter$count = 1748;
	#10 counter$count = 1749;
	#10 counter$count = 1750;
	#10 counter$count = 1751;
	#10 counter$count = 1752;
	#10 counter$count = 1753;
	#10 counter$count = 1754;
	#10 counter$count = 1755;
	#10 counter$count = 1756;
	#10 counter$count = 1757;
	#10 counter$count = 1758;
	#10 counter$count = 1759;
	#10 counter$count = 1760;
	#10 counter$count = 1761;
	#10 counter$count = 1762;
	#10 counter$count = 1763;
	#10 counter$count = 1764;
	#10 counter$count = 1765;
	#10 counter$count = 1766;
	#10 counter$count = 1767;
	#10 counter$count = 1768;
	#10 counter$count = 1769;
	#10 counter$count = 1770;
	#10 counter$count = 1771;
	#10 counter$count = 1772;
	#10 counter$count = 1773;
	#10 counter$count = 1774;
	#10 counter$count = 1775;
	#10 counter$count = 1776;
	#10 counter$count = 1777;
	#10 counter$count = 1778;
	#10 counter$count = 1779;
	#10 counter$count = 1780;
	#10 counter$count = 1781;
	#10 counter$count = 1782;
	#10 counter$count = 1783;
	#10 counter$count = 1784;
	#10 counter$count = 1785;
	#10 counter$count = 1786;
	#10 counter$count = 1787;
	#10 counter$count = 1788;
	#10 counter$count = 1789;
	#10 counter$count = 1790;
	#10 counter$count = 1791;
	#10 counter$count = 1792;
	#10 counter$count = 1793;
	#10 counter$count = 1794;
	#10 counter$count = 1795;
	#10 counter$count = 1796;
	#10 counter$count = 1797;
	#10 counter$count = 1798;
	#10 counter$count = 1799;
	#10 counter$count = 1800;
	#10 counter$count = 1801;
	#10 counter$count = 1802;
	#10 counter$count = 1803;
	#10 counter$count = 1804;
	#10 counter$count = 1805;
	#10 counter$count = 1806;
	#10 counter$count = 1807;
	#10 counter$count = 1808;
	#10 counter$count = 1809;
	#10 counter$count = 1810;
	#10 counter$count = 1811;
	#10 counter$count = 1812;
	#10 counter$count = 1813;
	#10 counter$count = 1814;
	#10 counter$count = 1815;
	#10 counter$count = 1816;
	#10 counter$count = 1817;
	#10 counter$count = 1818;
	#10 counter$count = 1819;
	#10 counter$count = 1820;
	#10 counter$count = 1821;
	#10 counter$count = 1822;
	#10 counter$count = 1823;
	#10 counter$count = 1824;
	#10 counter$count = 1825;
	#10 counter$count = 1826;
	#10 counter$count = 1827;
	#10 counter$count = 1828;
	#10 counter$count = 1829;
	#10 counter$count = 1830;
	#10 counter$count = 1831;
	#10 counter$count = 1832;
	#10 counter$count = 1833;
	#10 counter$count = 1834;
	#10 counter$count = 1835;
	#10 counter$count = 1836;
	#10 counter$count = 1837;
	#10 counter$count = 1838;
	#10 counter$count = 1839;
	#10 counter$count = 1840;
	#10 counter$count = 1841;
	#10 counter$count = 1842;
	#10 counter$count = 1843;
	#10 counter$count = 1844;
	#10 counter$count = 1845;
	#10 counter$count = 1846;
	#10 counter$count = 1847;
	#10 counter$count = 1848;
	#10 counter$count = 1849;
	#10 counter$count = 1850;
	#10 counter$count = 1851;
	#10 counter$count = 1852;
	#10 counter$count = 1853;
	#10 counter$count = 1854;
	#10 counter$count = 1855;
	#10 counter$count = 1856;
	#10 counter$count = 1857;
	#10 counter$count = 1858;
	#10 counter$count = 1859;
	#10 counter$count = 1860;
	#10 counter$count = 1861;
	#10 counter$count = 1862;
	#10 counter$count = 1863;
	#10 counter$count = 1864;
	#10 counter$count = 1865;
	#10 counter$count = 1866;
	#10 counter$count = 1867;
	#10 counter$count = 1868;
	#10 counter$count = 1869;
	#10 counter$count = 1870;
	#10 counter$count = 1871;
	#10 counter$count = 1872;
	#10 counter$count = 1873;
	#10 counter$count = 1874;
	#10 counter$count = 1875;
	#10 counter$count = 1876;
	#10 counter$count = 1877;
	#10 counter$count = 1878;
	#10 counter$count = 1879;
	#10 counter$count = 1880;
	#10 counter$count = 1881;
	#10 counter$count = 1882;
	#10 counter$count = 1883;
	#10 counter$count = 1884;
	#10 counter$count = 1885;
	#10 counter$count = 1886;
	#10 counter$count = 1887;
	#10 counter$count = 1888;
	#10 counter$count = 1889;
	#10 counter$count = 1890;
	#10 counter$count = 1891;
	#10 counter$count = 1892;
	#10 counter$count = 1893;
	#10 counter$count = 1894;
	#10 counter$count = 1895;
	#10 counter$count = 1896;
	#10 counter$count = 1897;
	#10 counter$count = 1898;
	#10 counter$count = 1899;
	#10 counter$count = 1900;
	#10 counter$count = 1901;
	#10 counter$count = 1902;
	#10 counter$count = 1903;
	#10 counter$count = 1904;
	#10 counter$count = 1905;
	#10 counter$count = 1906;
	#10 counter$count = 1907;
	#10 counter$count = 1908;
	#10 counter$count = 1909;
	#10 counter$count = 1910;
	#10 counter$count = 1911;
	#10 counter$count = 1912;
	#10 counter$count = 1913;
	#10 counter$count = 1914;
	#10 counter$count = 1915;
	#10 counter$count = 1916;
	#10 counter$count = 1917;
	#10 counter$count = 1918;
	#10 counter$count = 1919;
	#10 counter$count = 1920;
	#10 counter$count = 1921;
	#10 counter$count = 1922;
	#10 counter$count = 1923;
	#10 counter$count = 1924;
	#10 counter$count = 1925;
	#10 counter$count = 1926;
	#10 counter$count = 1927;
	#10 counter$count = 1928;
	#10 counter$count = 1929;
	#10 counter$count = 1930;
	#10 counter$count = 1931;
	#10 counter$count = 1932;
	#10 counter$count = 1933;
	#10 counter$count = 1934;
	#10 counter$count = 1935;
	#10 counter$count = 1936;
	#10 counter$count = 1937;
	#10 counter$count = 1938;
	#10 counter$count = 1939;
	#10 counter$count = 1940;
	#10 counter$count = 1941;
	#10 counter$count = 1942;
	#10 counter$count = 1943;
	#10 counter$count = 1944;
	#10 counter$count = 1945;
	#10 counter$count = 1946;
	#10 counter$count = 1947;
	#10 counter$count = 1948;
	#10 counter$count = 1949;
	#10 counter$count = 1950;
	#10 counter$count = 1951;
	#10 counter$count = 1952;
	#10 counter$count = 1953;
	#10 counter$count = 1954;
	#10 counter$count = 1955;
	#10 counter$count = 1956;
	#10 counter$count = 1957;
	#10 counter$count = 1958;
	#10 counter$count = 1959;
	#10 counter$count = 1960;
	#10 counter$count = 1961;
	#10 counter$count = 1962;
	#10 counter$count = 1963;
	#10 counter$count = 1964;
	#10 counter$count = 1965;
	#10 counter$count = 1966;
	#10 counter$count = 1967;
	#10 counter$count = 1968;
	#10 counter$count = 1969;
	#10 counter$count = 1970;
	#10 counter$count = 1971;
	#10 counter$count = 1972;
	#10 counter$count = 1973;
	#10 counter$count = 1974;
	#10 counter$count = 1975;
	#10 counter$count = 1976;
	#10 counter$count = 1977;
	#10 counter$count = 1978;
	#10 counter$count = 1979;
	#10 counter$count = 1980;
	#10 counter$count = 1981;
	#10 counter$count = 1982;
	#10 counter$count = 1983;
	#10 counter$count = 1984;
	#10 counter$count = 1985;
	#10 counter$count = 1986;
	#10 counter$count = 1987;
	#10 counter$count = 1988;
	#10 counter$count = 1989;
	#10 counter$count = 1990;
	#10 counter$count = 1991;
	#10 counter$count = 1992;
	#10 counter$count = 1993;
	#10 counter$count = 1994;
	#10 counter$count = 1995;
	#10 counter$count = 1996;
	#10 counter$count = 1997;
	#10 counter$count = 1998;
	#10 counter$count = 1999;
	#10 counter$count = 2000;
	#10 counter$count = 2001;
	#10 counter$count = 2002;
	#10 counter$count = 2003;
	#10 counter$count = 2004;
	#10 counter$count = 2005;
	#10 counter$count = 2006;
	#10 counter$count = 2007;
	#10 counter$count = 2008;
	#10 counter$count = 2009;
	#10 counter$count = 2010;
	#10 counter$count = 2011;
	#10 counter$count = 2012;
	#10 counter$count = 2013;
	#10 counter$count = 2014;
	#10 counter$count = 2015;
	#10 counter$count = 2016;
	#10 counter$count = 2017;
	#10 counter$count = 2018;
	#10 counter$count = 2019;
	#10 counter$count = 2020;
	#10 counter$count = 2021;
	#10 counter$count = 2022;
	#10 counter$count = 2023;
	#10 counter$count = 2024;
	#10 counter$count = 2025;
	#10 counter$count = 2026;
	#10 counter$count = 2027;
	#10 counter$count = 2028;
	#10 counter$count = 2029;
	#10 counter$count = 2030;
	#10 counter$count = 2031;
	#10 counter$count = 2032;
	#10 counter$count = 2033;
	#10 counter$count = 2034;
	#10 counter$count = 2035;
	#10 counter$count = 2036;
	#10 counter$count = 2037;
	#10 counter$count = 2038;
	#10 counter$count = 2039;
	#10 counter$count = 2040;
	#10 counter$count = 2041;
	#10 counter$count = 2042;
	#10 counter$count = 2043;
	#10 counter$count = 2044;
	#10 counter$count = 2045;
	#10 counter$count = 2046;
	#10 counter$count = 2047;
	#10 counter$count = 2048;
	#10 counter$count = 2049;
	#10 counter$count = 2050;
	#10 counter$count = 2051;
	#10 counter$count = 2052;
	#10 counter$count = 2053;
	#10 counter$count = 2054;
	#10 counter$count = 2055;
	#10 counter$count = 2056;
	#10 counter$count = 2057;
	#10 counter$count = 2058;
	#10 counter$count = 2059;
	#10 counter$count = 2060;
	#10 counter$count = 2061;
	#10 counter$count = 2062;
	#10 counter$count = 2063;
	#10 counter$count = 2064;
	#10 counter$count = 2065;
	#10 counter$count = 2066;
	#10 counter$count = 2067;
	#10 counter$count = 2068;
	#10 counter$count = 2069;
	#10 counter$count = 2070;
	#10 counter$count = 2071;
	#10 counter$count = 2072;
	#10 counter$count = 2073;
	#10 counter$count = 2074;
	#10 counter$count = 2075;
	#10 counter$count = 2076;
	#10 counter$count = 2077;
	#10 counter$count = 2078;
	#10 counter$count = 2079;
	#10 counter$count = 2080;
	#10 counter$count = 2081;
	#10 counter$count = 2082;
	#10 counter$count = 2083;
	#10 counter$count = 2084;
	#10 counter$count = 2085;
	#10 counter$count = 2086;
	#10 counter$count = 2087;
	#10 counter$count = 2088;
	#10 counter$count = 2089;
	#10 counter$count = 2090;
	#10 counter$count = 2091;
	#10 counter$count = 2092;
	#10 counter$count = 2093;
	#10 counter$count = 2094;
	#10 counter$count = 2095;
	#10 counter$count = 2096;
	#10 counter$count = 2097;
	#10 counter$count = 2098;
	#10 counter$count = 2099;
	#10 counter$count = 2100;
	#10 counter$count = 2101;
	#10 counter$count = 2102;
	#10 counter$count = 2103;
	#10 counter$count = 2104;
	#10 counter$count = 2105;
	#10 counter$count = 2106;
	#10 counter$count = 2107;
	#10 counter$count = 2108;
	#10 counter$count = 2109;
	#10 counter$count = 2110;
	#10 counter$count = 2111;
	#10 counter$count = 2112;
	#10 counter$count = 2113;
	#10 counter$count = 2114;
	#10 counter$count = 2115;
	#10 counter$count = 2116;
	#10 counter$count = 2117;
	#10 counter$count = 2118;
	#10 counter$count = 2119;
	#10 counter$count = 2120;
	#10 counter$count = 2121;
	#10 counter$count = 2122;
	#10 counter$count = 2123;
	#10 counter$count = 2124;
	#10 counter$count = 2125;
	#10 counter$count = 2126;
	#10 counter$count = 2127;
	#10 counter$count = 2128;
	#10 counter$count = 2129;
	#10 counter$count = 2130;
	#10 counter$count = 2131;
	#10 counter$count = 2132;
	#10 counter$count = 2133;
	#10 counter$count = 2134;
	#10 counter$count = 2135;
	#10 counter$count = 2136;
	#10 counter$count = 2137;
	#10 counter$count = 2138;
	#10 counter$count = 2139;
	#10 counter$count = 2140;
	#10 counter$count = 2141;
	#10 counter$count = 2142;
	#10 counter$count = 2143;
	#10 counter$count = 2144;
	#10 counter$count = 2145;
	#10 counter$count = 2146;
	#10 counter$count = 2147;
	#10 counter$count = 2148;
	#10 counter$count = 2149;
	#10 counter$count = 2150;
	#10 counter$count = 2151;
	#10 counter$count = 2152;
	#10 counter$count = 2153;
	#10 counter$count = 2154;
	#10 counter$count = 2155;
	#10 counter$count = 2156;
	#10 counter$count = 2157;
	#10 counter$count = 2158;
	#10 counter$count = 2159;
	#10 counter$count = 2160;
	#10 counter$count = 2161;
	#10 counter$count = 2162;
	#10 counter$count = 2163;
	#10 counter$count = 2164;
	#10 counter$count = 2165;
	#10 counter$count = 2166;
	#10 counter$count = 2167;
	#10 counter$count = 2168;
	#10 counter$count = 2169;
	#10 counter$count = 2170;
	#10 counter$count = 2171;
	#10 counter$count = 2172;
	#10 counter$count = 2173;
	#10 counter$count = 2174;
	#10 counter$count = 2175;
	#10 counter$count = 2176;
	#10 counter$count = 2177;
	#10 counter$count = 2178;
	#10 counter$count = 2179;
	#10 counter$count = 2180;
	#10 counter$count = 2181;
	#10 counter$count = 2182;
	#10 counter$count = 2183;
	#10 counter$count = 2184;
	#10 counter$count = 2185;
	#10 counter$count = 2186;
	#10 counter$count = 2187;
	#10 counter$count = 2188;
	#10 counter$count = 2189;
	#10 counter$count = 2190;
	#10 counter$count = 2191;
	#10 counter$count = 2192;
	#10 counter$count = 2193;
	#10 counter$count = 2194;
	#10 counter$count = 2195;
	#10 counter$count = 2196;
	#10 counter$count = 2197;
	#10 counter$count = 2198;
	#10 counter$count = 2199;
	#10 counter$count = 2200;
	#10 counter$count = 2201;
	#10 counter$count = 2202;
	#10 counter$count = 2203;
	#10 counter$count = 2204;
	#10 counter$count = 2205;
	#10 counter$count = 2206;
	#10 counter$count = 2207;
	#10 counter$count = 2208;
	#10 counter$count = 2209;
	#10 counter$count = 2210;
	#10 counter$count = 2211;
	#10 counter$count = 2212;
	#10 counter$count = 2213;
	#10 counter$count = 2214;
	#10 counter$count = 2215;
	#10 counter$count = 2216;
	#10 counter$count = 2217;
	#10 counter$count = 2218;
	#10 counter$count = 2219;
	#10 counter$count = 2220;
	#10 counter$count = 2221;
	#10 counter$count = 2222;
	#10 counter$count = 2223;
	#10 counter$count = 2224;
	#10 counter$count = 2225;
	#10 counter$count = 2226;
	#10 counter$count = 2227;
	#10 counter$count = 2228;
	#10 counter$count = 2229;
	#10 counter$count = 2230;
	#10 counter$count = 2231;
	#10 counter$count = 2232;
	#10 counter$count = 2233;
	#10 counter$count = 2234;
	#10 counter$count = 2235;
	#10 counter$count = 2236;
	#10 counter$count = 2237;
	#10 counter$count = 2238;
	#10 counter$count = 2239;
	#10 counter$count = 2240;
	#10 counter$count = 2241;
	#10 counter$count = 2242;
	#10 counter$count = 2243;
	#10 counter$count = 2244;
	#10 counter$count = 2245;
	#10 counter$count = 2246;
	#10 counter$count = 2247;
	#10 counter$count = 2248;
	#10 counter$count = 2249;
	#10 counter$count = 2250;
	#10 counter$count = 2251;
	#10 counter$count = 2252;
	#10 counter$count = 2253;
	#10 counter$count = 2254;
	#10 counter$count = 2255;
	#10 counter$count = 2256;
	#10 counter$count = 2257;
	#10 counter$count = 2258;
	#10 counter$count = 2259;
	#10 counter$count = 2260;
	#10 counter$count = 2261;
	#10 counter$count = 2262;
	#10 counter$count = 2263;
	#10 counter$count = 2264;
	#10 counter$count = 2265;
	#10 counter$count = 2266;
	#10 counter$count = 2267;
	#10 counter$count = 2268;
	#10 counter$count = 2269;
	#10 counter$count = 2270;
	#10 counter$count = 2271;
	#10 counter$count = 2272;
	#10 counter$count = 2273;
	#10 counter$count = 2274;
	#10 counter$count = 2275;
	#10 counter$count = 2276;
	#10 counter$count = 2277;
	#10 counter$count = 2278;
	#10 counter$count = 2279;
	#10 counter$count = 2280;
	#10 counter$count = 2281;
	#10 counter$count = 2282;
	#10 counter$count = 2283;
	#10 counter$count = 2284;
	#10 counter$count = 2285;
	#10 counter$count = 2286;
	#10 counter$count = 2287;
	#10 counter$count = 2288;
	#10 counter$count = 2289;
	#10 counter$count = 2290;
	#10 counter$count = 2291;
	#10 counter$count = 2292;
	#10 counter$count = 2293;
	#10 counter$count = 2294;
	#10 counter$count = 2295;
	#10 counter$count = 2296;
	#10 counter$count = 2297;
	#10 counter$count = 2298;
	#10 counter$count = 2299;
	#10 counter$count = 2300;
	#10 counter$count = 2301;
	#10 counter$count = 2302;
	#10 counter$count = 2303;
	#10 counter$count = 2304;
	#10 counter$count = 2305;
	#10 counter$count = 2306;
	#10 counter$count = 2307;
	#10 counter$count = 2308;
	#10 counter$count = 2309;
	#10 counter$count = 2310;
	#10 counter$count = 2311;
	#10 counter$count = 2312;
	#10 counter$count = 2313;
	#10 counter$count = 2314;
	#10 counter$count = 2315;
	#10 counter$count = 2316;
	#10 counter$count = 2317;
	#10 counter$count = 2318;
	#10 counter$count = 2319;
	#10 counter$count = 2320;
	#10 counter$count = 2321;
	#10 counter$count = 2322;
	#10 counter$count = 2323;
	#10 counter$count = 2324;
	#10 counter$count = 2325;
	#10 counter$count = 2326;
	#10 counter$count = 2327;
	#10 counter$count = 2328;
	#10 counter$count = 2329;
	#10 counter$count = 2330;
	#10 counter$count = 2331;
	#10 counter$count = 2332;
	#10 counter$count = 2333;
	#10 counter$count = 2334;
	#10 counter$count = 2335;
	#10 counter$count = 2336;
	#10 counter$count = 2337;
	#10 counter$count = 2338;
	#10 counter$count = 2339;
	#10 counter$count = 2340;
	#10 counter$count = 2341;
	#10 counter$count = 2342;
	#10 counter$count = 2343;
	#10 counter$count = 2344;
	#10 counter$count = 2345;
	#10 counter$count = 2346;
	#10 counter$count = 2347;
	#10 counter$count = 2348;
	#10 counter$count = 2349;
	#10 counter$count = 2350;
	#10 counter$count = 2351;
	#10 counter$count = 2352;
	#10 counter$count = 2353;
	#10 counter$count = 2354;
	#10 counter$count = 2355;
	#10 counter$count = 2356;
	#10 counter$count = 2357;
	#10 counter$count = 2358;
	#10 counter$count = 2359;
	#10 counter$count = 2360;
	#10 counter$count = 2361;
	#10 counter$count = 2362;
	#10 counter$count = 2363;
	#10 counter$count = 2364;
	#10 counter$count = 2365;
	#10 counter$count = 2366;
	#10 counter$count = 2367;
	#10 counter$count = 2368;
	#10 counter$count = 2369;
	#10 counter$count = 2370;
	#10 counter$count = 2371;
	#10 counter$count = 2372;
	#10 counter$count = 2373;
	#10 counter$count = 2374;
	#10 counter$count = 2375;
	#10 counter$count = 2376;
	#10 counter$count = 2377;
	#10 counter$count = 2378;
	#10 counter$count = 2379;
	#10 counter$count = 2380;
	#10 counter$count = 2381;
	#10 counter$count = 2382;
	#10 counter$count = 2383;
	#10 counter$count = 2384;
	#10 counter$count = 2385;
	#10 counter$count = 2386;
	#10 counter$count = 2387;
	#10 counter$count = 2388;
	#10 counter$count = 2389;
	#10 counter$count = 2390;
	#10 counter$count = 2391;
	#10 counter$count = 2392;
	#10 counter$count = 2393;
	#10 counter$count = 2394;
	#10 counter$count = 2395;
	#10 counter$count = 2396;
	#10 counter$count = 2397;
	#10 counter$count = 2398;
	#10 counter$count = 2399;
	#10 counter$count = 2400;
	#10 counter$count = 2401;
	#10 counter$count = 2402;
	#10 counter$count = 2403;
	#10 counter$count = 2404;
	#10 counter$count = 2405;
	#10 counter$count = 2406;
	#10 counter$count = 2407;
	#10 counter$count = 2408;
	#10 counter$count = 2409;
	#10 counter$count = 2410;
	#10 counter$count = 2411;
	#10 counter$count = 2412;
	#10 counter$count = 2413;
	#10 counter$count = 2414;
	#10 counter$count = 2415;
	#10 counter$count = 2416;
	#10 counter$count = 2417;
	#10 counter$count = 2418;
	#10 counter$count = 2419;
	#10 counter$count = 2420;
	#10 counter$count = 2421;
	#10 counter$count = 2422;
	#10 counter$count = 2423;
	#10 counter$count = 2424;
	#10 counter$count = 2425;
	#10 counter$count = 2426;
	#10 counter$count = 2427;
	#10 counter$count = 2428;
	#10 counter$count = 2429;
	#10 counter$count = 2430;
	#10 counter$count = 2431;
	#10 counter$count = 2432;
	#10 counter$count = 2433;
	#10 counter$count = 2434;
	#10 counter$count = 2435;
	#10 counter$count = 2436;
	#10 counter$count = 2437;
	#10 counter$count = 2438;
	#10 counter$count = 2439;
	#10 counter$count = 2440;
	#10 counter$count = 2441;
	#10 counter$count = 2442;
	#10 counter$count = 2443;
	#10 counter$count = 2444;
	#10 counter$count = 2445;
	#10 counter$count = 2446;
	#10 counter$count = 2447;
	#10 counter$count = 2448;
	#10 counter$count = 2449;
	#10 counter$count = 2450;
	#10 counter$count = 2451;
	#10 counter$count = 2452;
	#10 counter$count = 2453;
	#10 counter$count = 2454;
	#10 counter$count = 2455;
	#10 counter$count = 2456;
	#10 counter$count = 2457;
	#10 counter$count = 2458;
	#10 counter$count = 2459;
	#10 counter$count = 2460;
	#10 counter$count = 2461;
	#10 counter$count = 2462;
	#10 counter$count = 2463;
	#10 counter$count = 2464;
	#10 counter$count = 2465;
	#10 counter$count = 2466;
	#10 counter$count = 2467;
	#10 counter$count = 2468;
	#10 counter$count = 2469;
	#10 counter$count = 2470;
	#10 counter$count = 2471;
	#10 counter$count = 2472;
	#10 counter$count = 2473;
	#10 counter$count = 2474;
	#10 counter$count = 2475;
	#10 counter$count = 2476;
	#10 counter$count = 2477;
	#10 counter$count = 2478;
	#10 counter$count = 2479;
	#10 counter$count = 2480;
	#10 counter$count = 2481;
	#10 counter$count = 2482;
	#10 counter$count = 2483;
	#10 counter$count = 2484;
	#10 counter$count = 2485;
	#10 counter$count = 2486;
	#10 counter$count = 2487;
	#10 counter$count = 2488;
	#10 counter$count = 2489;
	#10 counter$count = 2490;
	#10 counter$count = 2491;
	#10 counter$count = 2492;
	#10 counter$count = 2493;
	#10 counter$count = 2494;
	#10 counter$count = 2495;
	#10 counter$count = 2496;
	#10 counter$count = 2497;
	#10 counter$count = 2498;
	#10 counter$count = 2499;
	#10 counter$count = 2500;
	#10 counter$count = 2501;
	#10 counter$count = 2502;
	#10 counter$count = 2503;
	#10 counter$count = 2504;
	#10 counter$count = 2505;
	#10 counter$count = 2506;
	#10 counter$count = 2507;
	#10 counter$count = 2508;
	#10 counter$count = 2509;
	#10 counter$count = 2510;
	#10 counter$count = 2511;
	#10 counter$count = 2512;
	#10 counter$count = 2513;
	#10 counter$count = 2514;
	#10 counter$count = 2515;
	#10 counter$count = 2516;
	#10 counter$count = 2517;
	#10 counter$count = 2518;
	#10 counter$count = 2519;
	#10 counter$count = 2520;
	#10 counter$count = 2521;
	#10 counter$count = 2522;
	#10 counter$count = 2523;
	#10 counter$count = 2524;
	#10 counter$count = 2525;
	#10 counter$count = 2526;
	#10 counter$count = 2527;
	#10 counter$count = 2528;
	#10 counter$count = 2529;
	#10 counter$count = 2530;
	#10 counter$count = 2531;
	#10 counter$count = 2532;
	#10 counter$count = 2533;
	#10 counter$count = 2534;
	#10 counter$count = 2535;
	#10 counter$count = 2536;
	#10 counter$count = 2537;
	#10 counter$count = 2538;
	#10 counter$count = 2539;
	#10 counter$count = 2540;
	#10 counter$count = 2541;
	#10 counter$count = 2542;
	#10 counter$count = 2543;
	#10 counter$count = 2544;
	#10 counter$count = 2545;
	#10 counter$count = 2546;
	#10 counter$count = 2547;
	#10 counter$count = 2548;
	#10 counter$count = 2549;
	#10 counter$count = 2550;
	#10 counter$count = 2551;
	#10 counter$count = 2552;
	#10 counter$count = 2553;
	#10 counter$count = 2554;
	#10 counter$count = 2555;
	#10 counter$count = 2556;
	#10 counter$count = 2557;
	#10 counter$count = 2558;
	#10 counter$count = 2559;
	#10 counter$count = 2560;
	#10 counter$count = 2561;
	#10 counter$count = 2562;
	#10 counter$count = 2563;
	#10 counter$count = 2564;
	#10 counter$count = 2565;
	#10 counter$count = 2566;
	#10 counter$count = 2567;
	#10 counter$count = 2568;
	#10 counter$count = 2569;
	#10 counter$count = 2570;
	#10 counter$count = 2571;
	#10 counter$count = 2572;
	#10 counter$count = 2573;
	#10 counter$count = 2574;
	#10 counter$count = 2575;
	#10 counter$count = 2576;
	#10 counter$count = 2577;
	#10 counter$count = 2578;
	#10 counter$count = 2579;
	#10 counter$count = 2580;
	#10 counter$count = 2581;
	#10 counter$count = 2582;
	#10 counter$count = 2583;
	#10 counter$count = 2584;
	#10 counter$count = 2585;
	#10 counter$count = 2586;
	#10 counter$count = 2587;
	#10 counter$count = 2588;
	#10 counter$count = 2589;
	#10 counter$count = 2590;
	#10 counter$count = 2591;
	#10 counter$count = 2592;
	#10 counter$count = 2593;
	#10 counter$count = 2594;
	#10 counter$count = 2595;
	#10 counter$count = 2596;
	#10 counter$count = 2597;
	#10 counter$count = 2598;
	#10 counter$count = 2599;
	#10 counter$count = 2600;
	#10 counter$count = 2601;
	#10 counter$count = 2602;
	#10 counter$count = 2603;
	#10 counter$count = 2604;
	#10 counter$count = 2605;
	#10 counter$count = 2606;
	#10 counter$count = 2607;
	#10 counter$count = 2608;
	#10 counter$count = 2609;
	#10 counter$count = 2610;
	#10 counter$count = 2611;
	#10 counter$count = 2612;
	#10 counter$count = 2613;
	#10 counter$count = 2614;
	#10 counter$count = 2615;
	#10 counter$count = 2616;
	#10 counter$count = 2617;
	#10 counter$count = 2618;
	#10 counter$count = 2619;
	#10 counter$count = 2620;
	#10 counter$count = 2621;
	#10 counter$count = 2622;
	#10 counter$count = 2623;
	#10 counter$count = 2624;
	#10 counter$count = 2625;
	#10 counter$count = 2626;
	#10 counter$count = 2627;
	#10 counter$count = 2628;
	#10 counter$count = 2629;
	#10 counter$count = 2630;
	#10 counter$count = 2631;
	#10 counter$count = 2632;
	#10 counter$count = 2633;
	#10 counter$count = 2634;
	#10 counter$count = 2635;
	#10 counter$count = 2636;
	#10 counter$count = 2637;
	#10 counter$count = 2638;
	#10 counter$count = 2639;
	#10 counter$count = 2640;
	#10 counter$count = 2641;
	#10 counter$count = 2642;
	#10 counter$count = 2643;
	#10 counter$count = 2644;
	#10 counter$count = 2645;
	#10 counter$count = 2646;
	#10 counter$count = 2647;
	#10 counter$count = 2648;
	#10 counter$count = 2649;
	#10 counter$count = 2650;
	#10 counter$count = 2651;
	#10 counter$count = 2652;
	#10 counter$count = 2653;
	#10 counter$count = 2654;
	#10 counter$count = 2655;
	#10 counter$count = 2656;
	#10 counter$count = 2657;
	#10 counter$count = 2658;
	#10 counter$count = 2659;
	#10 counter$count = 2660;
	#10 counter$count = 2661;
	#10 counter$count = 2662;
	#10 counter$count = 2663;
	#10 counter$count = 2664;
	#10 counter$count = 2665;
	#10 counter$count = 2666;
	#10 counter$count = 2667;
	#10 counter$count = 2668;
	#10 counter$count = 2669;
	#10 counter$count = 2670;
	#10 counter$count = 2671;
	#10 counter$count = 2672;
	#10 counter$count = 2673;
	#10 counter$count = 2674;
	#10 counter$count = 2675;
	#10 counter$count = 2676;
	#10 counter$count = 2677;
	#10 counter$count = 2678;
	#10 counter$count = 2679;
	#10 counter$count = 2680;
	#10 counter$count = 2681;
	#10 counter$count = 2682;
	#10 counter$count = 2683;
	#10 counter$count = 2684;
	#10 counter$count = 2685;
	#10 counter$count = 2686;
	#10 counter$count = 2687;
	#10 counter$count = 2688;
	#10 counter$count = 2689;
	#10 counter$count = 2690;
	#10 counter$count = 2691;
	#10 counter$count = 2692;
	#10 counter$count = 2693;
	#10 counter$count = 2694;
	#10 counter$count = 2695;
	#10 counter$count = 2696;
	#10 counter$count = 2697;
	#10 counter$count = 2698;
	#10 counter$count = 2699;
	#10 counter$count = 2700;
	#10 counter$count = 2701;
	#10 counter$count = 2702;
	#10 counter$count = 2703;
	#10 counter$count = 2704;
	#10 counter$count = 2705;
	#10 counter$count = 2706;
	#10 counter$count = 2707;
	#10 counter$count = 2708;
	#10 counter$count = 2709;
	#10 counter$count = 2710;
	#10 counter$count = 2711;
	#10 counter$count = 2712;
	#10 counter$count = 2713;
	#10 counter$count = 2714;
	#10 counter$count = 2715;
	#10 counter$count = 2716;
	#10 counter$count = 2717;
	#10 counter$count = 2718;
	#10 counter$count = 2719;
	#10 counter$count = 2720;
	#10 counter$count = 2721;
	#10 counter$count = 2722;
	#10 counter$count = 2723;
	#10 counter$count = 2724;
	#10 counter$count = 2725;
	#10 counter$count = 2726;
	#10 counter$count = 2727;
	#10 counter$count = 2728;
	#10 counter$count = 2729;
	#10 counter$count = 2730;
	#10 counter$count = 2731;
	#10 counter$count = 2732;
	#10 counter$count = 2733;
	#10 counter$count = 2734;
	#10 counter$count = 2735;
	#10 counter$count = 2736;
	#10 counter$count = 2737;
	#10 counter$count = 2738;
	#10 counter$count = 2739;
	#10 counter$count = 2740;
	#10 counter$count = 2741;
	#10 counter$count = 2742;
	#10 counter$count = 2743;
	#10 counter$count = 2744;
	#10 counter$count = 2745;
	#10 counter$count = 2746;
	#10 counter$count = 2747;
	#10 counter$count = 2748;
	#10 counter$count = 2749;
	#10 counter$count = 2750;
	#10 counter$count = 2751;
	#10 counter$count = 2752;
	#10 counter$count = 2753;
	#10 counter$count = 2754;
	#10 counter$count = 2755;
	#10 counter$count = 2756;
	#10 counter$count = 2757;
	#10 counter$count = 2758;
	#10 counter$count = 2759;
	#10 counter$count = 2760;
	#10 counter$count = 2761;
	#10 counter$count = 2762;
	#10 counter$count = 2763;
	#10 counter$count = 2764;
	#10 counter$count = 2765;
	#10 counter$count = 2766;
	#10 counter$count = 2767;
	#10 counter$count = 2768;
	#10 counter$count = 2769;
	#10 counter$count = 2770;
	#10 counter$count = 2771;
	#10 counter$count = 2772;
	#10 counter$count = 2773;
	#10 counter$count = 2774;
	#10 counter$count = 2775;
	#10 counter$count = 2776;
	#10 counter$count = 2777;
	#10 counter$count = 2778;
	#10 counter$count = 2779;
	#10 counter$count = 2780;
	#10 counter$count = 2781;
	#10 counter$count = 2782;
	#10 counter$count = 2783;
	#10 counter$count = 2784;
	#10 counter$count = 2785;
	#10 counter$count = 2786;
	#10 counter$count = 2787;
	#10 counter$count = 2788;
	#10 counter$count = 2789;
	#10 counter$count = 2790;
	#10 counter$count = 2791;
	#10 counter$count = 2792;
	#10 counter$count = 2793;
	#10 counter$count = 2794;
	#10 counter$count = 2795;
	#10 counter$count = 2796;
	#10 counter$count = 2797;
	#10 counter$count = 2798;
	#10 counter$count = 2799;
	#10 counter$count = 2800;
	#10 counter$count = 2801;
	#10 counter$count = 2802;
	#10 counter$count = 2803;
	#10 counter$count = 2804;
	#10 counter$count = 2805;
	#10 counter$count = 2806;
	#10 counter$count = 2807;
	#10 counter$count = 2808;
	#10 counter$count = 2809;
	#10 counter$count = 2810;
	#10 counter$count = 2811;
	#10 counter$count = 2812;
	#10 counter$count = 2813;
	#10 counter$count = 2814;
	#10 counter$count = 2815;
	#10 counter$count = 2816;
	#10 counter$count = 2817;
	#10 counter$count = 2818;
	#10 counter$count = 2819;
	#10 counter$count = 2820;
	#10 counter$count = 2821;
	#10 counter$count = 2822;
	#10 counter$count = 2823;
	#10 counter$count = 2824;
	#10 counter$count = 2825;
	#10 counter$count = 2826;
	#10 counter$count = 2827;
	#10 counter$count = 2828;
	#10 counter$count = 2829;
	#10 counter$count = 2830;
	#10 counter$count = 2831;
	#10 counter$count = 2832;
	#10 counter$count = 2833;
	#10 counter$count = 2834;
	#10 counter$count = 2835;
	#10 counter$count = 2836;
	#10 counter$count = 2837;
	#10 counter$count = 2838;
	#10 counter$count = 2839;
	#10 counter$count = 2840;
	#10 counter$count = 2841;
	#10 counter$count = 2842;
	#10 counter$count = 2843;
	#10 counter$count = 2844;
	#10 counter$count = 2845;
	#10 counter$count = 2846;
	#10 counter$count = 2847;
	#10 counter$count = 2848;
	#10 counter$count = 2849;
	#10 counter$count = 2850;
	#10 counter$count = 2851;
	#10 counter$count = 2852;
	#10 counter$count = 2853;
	#10 counter$count = 2854;
	#10 counter$count = 2855;
	#10 counter$count = 2856;
	#10 counter$count = 2857;
	#10 counter$count = 2858;
	#10 counter$count = 2859;
	#10 counter$count = 2860;
	#10 counter$count = 2861;
	#10 counter$count = 2862;
	#10 counter$count = 2863;
	#10 counter$count = 2864;
	#10 counter$count = 2865;
	#10 counter$count = 2866;
	#10 counter$count = 2867;
	#10 counter$count = 2868;
	#10 counter$count = 2869;
	#10 counter$count = 2870;
	#10 counter$count = 2871;
	#10 counter$count = 2872;
	#10 counter$count = 2873;
	#10 counter$count = 2874;
	#10 counter$count = 2875;
	#10 counter$count = 2876;
	#10 counter$count = 2877;
	#10 counter$count = 2878;
	#10 counter$count = 2879;
	#10 counter$count = 2880;
	#10 counter$count = 2881;
	#10 counter$count = 2882;
	#10 counter$count = 2883;
	#10 counter$count = 2884;
	#10 counter$count = 2885;
	#10 counter$count = 2886;
	#10 counter$count = 2887;
	#10 counter$count = 2888;
	#10 counter$count = 2889;
	#10 counter$count = 2890;
	#10 counter$count = 2891;
	#10 counter$count = 2892;
	#10 counter$count = 2893;
	#10 counter$count = 2894;
	#10 counter$count = 2895;
	#10 counter$count = 2896;
	#10 counter$count = 2897;
	#10 counter$count = 2898;
	#10 counter$count = 2899;
	#10 counter$count = 2900;
	#10 counter$count = 2901;
	#10 counter$count = 2902;
	#10 counter$count = 2903;
	#10 counter$count = 2904;
	#10 counter$count = 2905;
	#10 counter$count = 2906;
	#10 counter$count = 2907;
	#10 counter$count = 2908;
	#10 counter$count = 2909;
	#10 counter$count = 2910;
	#10 counter$count = 2911;
	#10 counter$count = 2912;
	#10 counter$count = 2913;
	#10 counter$count = 2914;
	#10 counter$count = 2915;
	#10 counter$count = 2916;
	#10 counter$count = 2917;
	#10 counter$count = 2918;
	#10 counter$count = 2919;
	#10 counter$count = 2920;
	#10 counter$count = 2921;
	#10 counter$count = 2922;
	#10 counter$count = 2923;
	#10 counter$count = 2924;
	#10 counter$count = 2925;
	#10 counter$count = 2926;
	#10 counter$count = 2927;
	#10 counter$count = 2928;
	#10 counter$count = 2929;
	#10 counter$count = 2930;
	#10 counter$count = 2931;
	#10 counter$count = 2932;
	#10 counter$count = 2933;
	#10 counter$count = 2934;
	#10 counter$count = 2935;
	#10 counter$count = 2936;
	#10 counter$count = 2937;
	#10 counter$count = 2938;
	#10 counter$count = 2939;
	#10 counter$count = 2940;
	#10 counter$count = 2941;
	#10 counter$count = 2942;
	#10 counter$count = 2943;
	#10 counter$count = 2944;
	#10 counter$count = 2945;
	#10 counter$count = 2946;
	#10 counter$count = 2947;
	#10 counter$count = 2948;
	#10 counter$count = 2949;
	#10 counter$count = 2950;
	#10 counter$count = 2951;
	#10 counter$count = 2952;
	#10 counter$count = 2953;
	#10 counter$count = 2954;
	#10 counter$count = 2955;
	#10 counter$count = 2956;
	#10 counter$count = 2957;
	#10 counter$count = 2958;
	#10 counter$count = 2959;
	#10 counter$count = 2960;
	#10 counter$count = 2961;
	#10 counter$count = 2962;
	#10 counter$count = 2963;
	#10 counter$count = 2964;
	#10 counter$count = 2965;
	#10 counter$count = 2966;
	#10 counter$count = 2967;
	#10 counter$count = 2968;
	#10 counter$count = 2969;
	#10 counter$count = 2970;
	#10 counter$count = 2971;
	#10 counter$count = 2972;
	#10 counter$count = 2973;
	#10 counter$count = 2974;
	#10 counter$count = 2975;
	#10 counter$count = 2976;
	#10 counter$count = 2977;
	#10 counter$count = 2978;
	#10 counter$count = 2979;
	#10 counter$count = 2980;
	#10 counter$count = 2981;
	#10 counter$count = 2982;
	#10 counter$count = 2983;
	#10 counter$count = 2984;
	#10 counter$count = 2985;
	#10 counter$count = 2986;
	#10 counter$count = 2987;
	#10 counter$count = 2988;
	#10 counter$count = 2989;
	#10 counter$count = 2990;
	#10 counter$count = 2991;
	#10 counter$count = 2992;
	#10 counter$count = 2993;
	#10 counter$count = 2994;
	#10 counter$count = 2995;
	#10 counter$count = 2996;
	#10 counter$count = 2997;
	#10 counter$count = 2998;
	#10 counter$count = 2999;
	#10 counter$count = 3000;
	#10 counter$count = 3001;
	#10 counter$count = 3002;
	#10 counter$count = 3003;
	#10 counter$count = 3004;
	#10 counter$count = 3005;
	#10 counter$count = 3006;
	#10 counter$count = 3007;
	#10 counter$count = 3008;
	#10 counter$count = 3009;
	#10 counter$count = 3010;
	#10 counter$count = 3011;
	#10 counter$count = 3012;
	#10 counter$count = 3013;
	#10 counter$count = 3014;
	#10 counter$count = 3015;
	#10 counter$count = 3016;
	#10 counter$count = 3017;
	#10 counter$count = 3018;
	#10 counter$count = 3019;
	#10 counter$count = 3020;
	#10 counter$count = 3021;
	#10 counter$count = 3022;
	#10 counter$count = 3023;
	#10 counter$count = 3024;
	#10 counter$count = 3025;
	#10 counter$count = 3026;
	#10 counter$count = 3027;
	#10 counter$count = 3028;
	#10 counter$count = 3029;
	#10 counter$count = 3030;
	#10 counter$count = 3031;
	#10 counter$count = 3032;
	#10 counter$count = 3033;
	#10 counter$count = 3034;
	#10 counter$count = 3035;
	#10 counter$count = 3036;
	#10 counter$count = 3037;
	#10 counter$count = 3038;
	#10 counter$count = 3039;
	#10 counter$count = 3040;
	#10 counter$count = 3041;
	#10 counter$count = 3042;
	#10 counter$count = 3043;
	#10 counter$count = 3044;
	#10 counter$count = 3045;
	#10 counter$count = 3046;
	#10 counter$count = 3047;
	#10 counter$count = 3048;
	#10 counter$count = 3049;
	#10 counter$count = 3050;
	#10 counter$count = 3051;
	#10 counter$count = 3052;
	#10 counter$count = 3053;
	#10 counter$count = 3054;
	#10 counter$count = 3055;
	#10 counter$count = 3056;
	#10 counter$count = 3057;
	#10 counter$count = 3058;
	#10 counter$count = 3059;
	#10 counter$count = 3060;
	#10 counter$count = 3061;
	#10 counter$count = 3062;
	#10 counter$count = 3063;
	#10 counter$count = 3064;
	#10 counter$count = 3065;
	#10 counter$count = 3066;
	#10 counter$count = 3067;
	#10 counter$count = 3068;
	#10 counter$count = 3069;
	#10 counter$count = 3070;
	#10 counter$count = 3071;
	#10 counter$count = 3072;
	#10 counter$count = 3073;
	#10 counter$count = 3074;
	#10 counter$count = 3075;
	#10 counter$count = 3076;
	#10 counter$count = 3077;
	#10 counter$count = 3078;
	#10 counter$count = 3079;
	#10 counter$count = 3080;
	#10 counter$count = 3081;
	#10 counter$count = 3082;
	#10 counter$count = 3083;
	#10 counter$count = 3084;
	#10 counter$count = 3085;
	#10 counter$count = 3086;
	#10 counter$count = 3087;
	#10 counter$count = 3088;
	#10 counter$count = 3089;
	#10 counter$count = 3090;
	#10 counter$count = 3091;
	#10 counter$count = 3092;
	#10 counter$count = 3093;
	#10 counter$count = 3094;
	#10 counter$count = 3095;
	#10 counter$count = 3096;
	#10 counter$count = 3097;
	#10 counter$count = 3098;
	#10 counter$count = 3099;
	#10 counter$count = 3100;
	#10 counter$count = 3101;
	#10 counter$count = 3102;
	#10 counter$count = 3103;
	#10 counter$count = 3104;
	#10 counter$count = 3105;
	#10 counter$count = 3106;
	#10 counter$count = 3107;
	#10 counter$count = 3108;
	#10 counter$count = 3109;
	#10 counter$count = 3110;
	#10 counter$count = 3111;
	#10 counter$count = 3112;
	#10 counter$count = 3113;
	#10 counter$count = 3114;
	#10 counter$count = 3115;
	#10 counter$count = 3116;
	#10 counter$count = 3117;
	#10 counter$count = 3118;
	#10 counter$count = 3119;
	#10 counter$count = 3120;
	#10 counter$count = 3121;
	#10 counter$count = 3122;
	#10 counter$count = 3123;
	#10 counter$count = 3124;
	#10 counter$count = 3125;
	#10 counter$count = 3126;
	#10 counter$count = 3127;
	#10 counter$count = 3128;
	#10 counter$count = 3129;
	#10 counter$count = 3130;
	#10 counter$count = 3131;
	#10 counter$count = 3132;
	#10 counter$count = 3133;
	#10 counter$count = 3134;
	#10 counter$count = 3135;
	#10 counter$count = 3136;
	#10 counter$count = 3137;
	#10 counter$count = 3138;
	#10 counter$count = 3139;
	#10 counter$count = 3140;
	#10 counter$count = 3141;
	#10 counter$count = 3142;
	#10 counter$count = 3143;
	#10 counter$count = 3144;
	#10 counter$count = 3145;
	#10 counter$count = 3146;
	#10 counter$count = 3147;
	#10 counter$count = 3148;
	#10 counter$count = 3149;
	#10 counter$count = 3150;
	#10 counter$count = 3151;
	#10 counter$count = 3152;
	#10 counter$count = 3153;
	#10 counter$count = 3154;
	#10 counter$count = 3155;
	#10 counter$count = 3156;
	#10 counter$count = 3157;
	#10 counter$count = 3158;
	#10 counter$count = 3159;
	#10 counter$count = 3160;
	#10 counter$count = 3161;
	#10 counter$count = 3162;
	#10 counter$count = 3163;
	#10 counter$count = 3164;
	#10 counter$count = 3165;
	#10 counter$count = 3166;
	#10 counter$count = 3167;
	#10 counter$count = 3168;
	#10 counter$count = 3169;
	#10 counter$count = 3170;
	#10 counter$count = 3171;
	#10 counter$count = 3172;
	#10 counter$count = 3173;
	#10 counter$count = 3174;
	#10 counter$count = 3175;
	#10 counter$count = 3176;
	#10 counter$count = 3177;
	#10 counter$count = 3178;
	#10 counter$count = 3179;
	#10 counter$count = 3180;
	#10 counter$count = 3181;
	#10 counter$count = 3182;
	#10 counter$count = 3183;
	#10 counter$count = 3184;
	#10 counter$count = 3185;
	#10 counter$count = 3186;
	#10 counter$count = 3187;
	#10 counter$count = 3188;
	#10 counter$count = 3189;
	#10 counter$count = 3190;
	#10 counter$count = 3191;
	#10 counter$count = 3192;
	#10 counter$count = 3193;
	#10 counter$count = 3194;
	#10 counter$count = 3195;
	#10 counter$count = 3196;
	#10 counter$count = 3197;
	#10 counter$count = 3198;
	#10 counter$count = 3199;
	#10 counter$count = 3200;
	#10 counter$count = 3201;
	#10 counter$count = 3202;
	#10 counter$count = 3203;
	#10 counter$count = 3204;
	#10 counter$count = 3205;
	#10 counter$count = 3206;
	#10 counter$count = 3207;
	#10 counter$count = 3208;
	#10 counter$count = 3209;
	#10 counter$count = 3210;
	#10 counter$count = 3211;
	#10 counter$count = 3212;
	#10 counter$count = 3213;
	#10 counter$count = 3214;
	#10 counter$count = 3215;
	#10 counter$count = 3216;
	#10 counter$count = 3217;
	#10 counter$count = 3218;
	#10 counter$count = 3219;
	#10 counter$count = 3220;
	#10 counter$count = 3221;
	#10 counter$count = 3222;
	#10 counter$count = 3223;
	#10 counter$count = 3224;
	#10 counter$count = 3225;
	#10 counter$count = 3226;
	#10 counter$count = 3227;
	#10 counter$count = 3228;
	#10 counter$count = 3229;
	#10 counter$count = 3230;
	#10 counter$count = 3231;
	#10 counter$count = 3232;
	#10 counter$count = 3233;
	#10 counter$count = 3234;
	#10 counter$count = 3235;
	#10 counter$count = 3236;
	#10 counter$count = 3237;
	#10 counter$count = 3238;
	#10 counter$count = 3239;
	#10 counter$count = 3240;
	#10 counter$count = 3241;
	#10 counter$count = 3242;
	#10 counter$count = 3243;
	#10 counter$count = 3244;
	#10 counter$count = 3245;
	#10 counter$count = 3246;
	#10 counter$count = 3247;
	#10 counter$count = 3248;
	#10 counter$count = 3249;
	#10 counter$count = 3250;
	#10 counter$count = 3251;
	#10 counter$count = 3252;
	#10 counter$count = 3253;
	#10 counter$count = 3254;
	#10 counter$count = 3255;
	#10 counter$count = 3256;
	#10 counter$count = 3257;
	#10 counter$count = 3258;
	#10 counter$count = 3259;
	#10 counter$count = 3260;
	#10 counter$count = 3261;
	#10 counter$count = 3262;
	#10 counter$count = 3263;
	#10 counter$count = 3264;
	#10 counter$count = 3265;
	#10 counter$count = 3266;
	#10 counter$count = 3267;
	#10 counter$count = 3268;
	#10 counter$count = 3269;
	#10 counter$count = 3270;
	#10 counter$count = 3271;
	#10 counter$count = 3272;
	#10 counter$count = 3273;
	#10 counter$count = 3274;
	#10 counter$count = 3275;
	#10 counter$count = 3276;
	#10 counter$count = 3277;
	#10 counter$count = 3278;
	#10 counter$count = 3279;
	#10 counter$count = 3280;
	#10 counter$count = 3281;
	#10 counter$count = 3282;
	#10 counter$count = 3283;
	#10 counter$count = 3284;
	#10 counter$count = 3285;
	#10 counter$count = 3286;
	#10 counter$count = 3287;
	#10 counter$count = 3288;
	#10 counter$count = 3289;
	#10 counter$count = 3290;
	#10 counter$count = 3291;
	#10 counter$count = 3292;
	#10 counter$count = 3293;
	#10 counter$count = 3294;
	#10 counter$count = 3295;
	#10 counter$count = 3296;
	#10 counter$count = 3297;
	#10 counter$count = 3298;
	#10 counter$count = 3299;
	#10 counter$count = 3300;
	#10 counter$count = 3301;
	#10 counter$count = 3302;
	#10 counter$count = 3303;
	#10 counter$count = 3304;
	#10 counter$count = 3305;
	#10 counter$count = 3306;
	#10 counter$count = 3307;
	#10 counter$count = 3308;
	#10 counter$count = 3309;
	#10 counter$count = 3310;
	#10 counter$count = 3311;
	#10 counter$count = 3312;
	#10 counter$count = 3313;
	#10 counter$count = 3314;
	#10 counter$count = 3315;
	#10 counter$count = 3316;
	#10 counter$count = 3317;
	#10 counter$count = 3318;
	#10 counter$count = 3319;
	#10 counter$count = 3320;
	#10 counter$count = 3321;
	#10 counter$count = 3322;
	#10 counter$count = 3323;
	#10 counter$count = 3324;
	#10 counter$count = 3325;
	#10 counter$count = 3326;
	#10 counter$count = 3327;
	#10 counter$count = 3328;
	#10 counter$count = 3329;
	#10 counter$count = 3330;
	#10 counter$count = 3331;
	#10 counter$count = 3332;
	#10 counter$count = 3333;
	#10 counter$count = 3334;
	#10 counter$count = 3335;
	#10 counter$count = 3336;
	#10 counter$count = 3337;
	#10 counter$count = 3338;
	#10 counter$count = 3339;
	#10 counter$count = 3340;
	#10 counter$count = 3341;
	#10 counter$count = 3342;
	#10 counter$count = 3343;
	#10 counter$count = 3344;
	#10 counter$count = 3345;
	#10 counter$count = 3346;
	#10 counter$count = 3347;
	#10 counter$count = 3348;
	#10 counter$count = 3349;
	#10 counter$count = 3350;
	#10 counter$count = 3351;
	#10 counter$count = 3352;
	#10 counter$count = 3353;
	#10 counter$count = 3354;
	#10 counter$count = 3355;
	#10 counter$count = 3356;
	#10 counter$count = 3357;
	#10 counter$count = 3358;
	#10 counter$count = 3359;
	#10 counter$count = 3360;
	#10 counter$count = 3361;
	#10 counter$count = 3362;
	#10 counter$count = 3363;
	#10 counter$count = 3364;
	#10 counter$count = 3365;
	#10 counter$count = 3366;
	#10 counter$count = 3367;
	#10 counter$count = 3368;
	#10 counter$count = 3369;
	#10 counter$count = 3370;
	#10 counter$count = 3371;
	#10 counter$count = 3372;
	#10 counter$count = 3373;
	#10 counter$count = 3374;
	#10 counter$count = 3375;
	#10 counter$count = 3376;
	#10 counter$count = 3377;
	#10 counter$count = 3378;
	#10 counter$count = 3379;
	#10 counter$count = 3380;
	#10 counter$count = 3381;
	#10 counter$count = 3382;
	#10 counter$count = 3383;
	#10 counter$count = 3384;
	#10 counter$count = 3385;
	#10 counter$count = 3386;
	#10 counter$count = 3387;
	#10 counter$count = 3388;
	#10 counter$count = 3389;
	#10 counter$count = 3390;
	#10 counter$count = 3391;
	#10 counter$count = 3392;
	#10 counter$count = 3393;
	#10 counter$count = 3394;
	#10 counter$count = 3395;
	#10 counter$count = 3396;
	#10 counter$count = 3397;
	#10 counter$count = 3398;
	#10 counter$count = 3399;
	#10 counter$count = 3400;
	#10 counter$count = 3401;
	#10 counter$count = 3402;
	#10 counter$count = 3403;
	#10 counter$count = 3404;
	#10 counter$count = 3405;
	#10 counter$count = 3406;
	#10 counter$count = 3407;
	#10 counter$count = 3408;
	#10 counter$count = 3409;
	#10 counter$count = 3410;
	#10 counter$count = 3411;
	#10 counter$count = 3412;
	#10 counter$count = 3413;
	#10 counter$count = 3414;
	#10 counter$count = 3415;
	#10 counter$count = 3416;
	#10 counter$count = 3417;
	#10 counter$count = 3418;
	#10 counter$count = 3419;
	#10 counter$count = 3420;
	#10 counter$count = 3421;
	#10 counter$count = 3422;
	#10 counter$count = 3423;
	#10 counter$count = 3424;
	#10 counter$count = 3425;
	#10 counter$count = 3426;
	#10 counter$count = 3427;
	#10 counter$count = 3428;
	#10 counter$count = 3429;
	#10 counter$count = 3430;
	#10 counter$count = 3431;
	#10 counter$count = 3432;
	#10 counter$count = 3433;
	#10 counter$count = 3434;
	#10 counter$count = 3435;
	#10 counter$count = 3436;
	#10 counter$count = 3437;
	#10 counter$count = 3438;
	#10 counter$count = 3439;
	#10 counter$count = 3440;
	#10 counter$count = 3441;
	#10 counter$count = 3442;
	#10 counter$count = 3443;
	#10 counter$count = 3444;
	#10 counter$count = 3445;
	#10 counter$count = 3446;
	#10 counter$count = 3447;
	#10 counter$count = 3448;
	#10 counter$count = 3449;
	#10 counter$count = 3450;
	#10 counter$count = 3451;
	#10 counter$count = 3452;
	#10 counter$count = 3453;
	#10 counter$count = 3454;
	#10 counter$count = 3455;
	#10 counter$count = 3456;
	#10 counter$count = 3457;
	#10 counter$count = 3458;
	#10 counter$count = 3459;
	#10 counter$count = 3460;
	#10 counter$count = 3461;
	#10 counter$count = 3462;
	#10 counter$count = 3463;
	#10 counter$count = 3464;
	#10 counter$count = 3465;
	#10 counter$count = 3466;
	#10 counter$count = 3467;
	#10 counter$count = 3468;
	#10 counter$count = 3469;
	#10 counter$count = 3470;
	#10 counter$count = 3471;
	#10 counter$count = 3472;
	#10 counter$count = 3473;
	#10 counter$count = 3474;
	#10 counter$count = 3475;
	#10 counter$count = 3476;
	#10 counter$count = 3477;
	#10 counter$count = 3478;
	#10 counter$count = 3479;
	#10 counter$count = 3480;
	#10 counter$count = 3481;
	#10 counter$count = 3482;
	#10 counter$count = 3483;
	#10 counter$count = 3484;
	#10 counter$count = 3485;
	#10 counter$count = 3486;
	#10 counter$count = 3487;
	#10 counter$count = 3488;
	#10 counter$count = 3489;
	#10 counter$count = 3490;
	#10 counter$count = 3491;
	#10 counter$count = 3492;
	#10 counter$count = 3493;
	#10 counter$count = 3494;
	#10 counter$count = 3495;
	#10 counter$count = 3496;
	#10 counter$count = 3497;
	#10 counter$count = 3498;
	#10 counter$count = 3499;
	#10 counter$count = 3500;
	#10 counter$count = 3501;
	#10 counter$count = 3502;
	#10 counter$count = 3503;
	#10 counter$count = 3504;
	#10 counter$count = 3505;
	#10 counter$count = 3506;
	#10 counter$count = 3507;
	#10 counter$count = 3508;
	#10 counter$count = 3509;
	#10 counter$count = 3510;
	#10 counter$count = 3511;
	#10 counter$count = 3512;
	#10 counter$count = 3513;
	#10 counter$count = 3514;
	#10 counter$count = 3515;
	#10 counter$count = 3516;
	#10 counter$count = 3517;
	#10 counter$count = 3518;
	#10 counter$count = 3519;
	#10 counter$count = 3520;
	#10 counter$count = 3521;
	#10 counter$count = 3522;
	#10 counter$count = 3523;
	#10 counter$count = 3524;
	#10 counter$count = 3525;
	#10 counter$count = 3526;
	#10 counter$count = 3527;
	#10 counter$count = 3528;
	#10 counter$count = 3529;
	#10 counter$count = 3530;
	#10 counter$count = 3531;
	#10 counter$count = 3532;
	#10 counter$count = 3533;
	#10 counter$count = 3534;
	#10 counter$count = 3535;
	#10 counter$count = 3536;
	#10 counter$count = 3537;
	#10 counter$count = 3538;
	#10 counter$count = 3539;
	#10 counter$count = 3540;
	#10 counter$count = 3541;
	#10 counter$count = 3542;
	#10 counter$count = 3543;
	#10 counter$count = 3544;
	#10 counter$count = 3545;
	#10 counter$count = 3546;
	#10 counter$count = 3547;
	#10 counter$count = 3548;
	#10 counter$count = 3549;
	#10 counter$count = 3550;
	#10 counter$count = 3551;
	#10 counter$count = 3552;
	#10 counter$count = 3553;
	#10 counter$count = 3554;
	#10 counter$count = 3555;
	#10 counter$count = 3556;
	#10 counter$count = 3557;
	#10 counter$count = 3558;
	#10 counter$count = 3559;
	#10 counter$count = 3560;
	#10 counter$count = 3561;
	#10 counter$count = 3562;
	#10 counter$count = 3563;
	#10 counter$count = 3564;
	#10 counter$count = 3565;
	#10 counter$count = 3566;
	#10 counter$count = 3567;
	#10 counter$count = 3568;
	#10 counter$count = 3569;
	#10 counter$count = 3570;
	#10 counter$count = 3571;
	#10 counter$count = 3572;
	#10 counter$count = 3573;
	#10 counter$count = 3574;
	#10 counter$count = 3575;
	#10 counter$count = 3576;
	#10 counter$count = 3577;
	#10 counter$count = 3578;
	#10 counter$count = 3579;
	#10 counter$count = 3580;
	#10 counter$count = 3581;
	#10 counter$count = 3582;
	#10 counter$count = 3583;
	#10 counter$count = 3584;
	#10 counter$count = 3585;
	#10 counter$count = 3586;
	#10 counter$count = 3587;
	#10 counter$count = 3588;
	#10 counter$count = 3589;
	#10 counter$count = 3590;
	#10 counter$count = 3591;
	#10 counter$count = 3592;
	#10 counter$count = 3593;
	#10 counter$count = 3594;
	#10 counter$count = 3595;
	#10 counter$count = 3596;
	#10 counter$count = 3597;
	#10 counter$count = 3598;
	#10 counter$count = 3599;
	#10 counter$count = 3600;
	#10 counter$count = 3601;
	#10 counter$count = 3602;
	#10 counter$count = 3603;
	#10 counter$count = 3604;
	#10 counter$count = 3605;
	#10 counter$count = 3606;
	#10 counter$count = 3607;
	#10 counter$count = 3608;
	#10 counter$count = 3609;
	#10 counter$count = 3610;
	#10 counter$count = 3611;
	#10 counter$count = 3612;
	#10 counter$count = 3613;
	#10 counter$count = 3614;
	#10 counter$count = 3615;
	#10 counter$count = 3616;
	#10 counter$count = 3617;
	#10 counter$count = 3618;
	#10 counter$count = 3619;
	#10 counter$count = 3620;
	#10 counter$count = 3621;
	#10 counter$count = 3622;
	#10 counter$count = 3623;
	#10 counter$count = 3624;
	#10 counter$count = 3625;
	#10 counter$count = 3626;
	#10 counter$count = 3627;
	#10 counter$count = 3628;
	#10 counter$count = 3629;
	#10 counter$count = 3630;
	#10 counter$count = 3631;
	#10 counter$count = 3632;
	#10 counter$count = 3633;
	#10 counter$count = 3634;
	#10 counter$count = 3635;
	#10 counter$count = 3636;
	#10 counter$count = 3637;
	#10 counter$count = 3638;
	#10 counter$count = 3639;
	#10 counter$count = 3640;
	#10 counter$count = 3641;
	#10 counter$count = 3642;
	#10 counter$count = 3643;
	#10 counter$count = 3644;
	#10 counter$count = 3645;
	#10 counter$count = 3646;
	#10 counter$count = 3647;
	#10 counter$count = 3648;
	#10 counter$count = 3649;
	#10 counter$count = 3650;
	#10 counter$count = 3651;
	#10 counter$count = 3652;
	#10 counter$count = 3653;
	#10 counter$count = 3654;
	#10 counter$count = 3655;
	#10 counter$count = 3656;
	#10 counter$count = 3657;
	#10 counter$count = 3658;
	#10 counter$count = 3659;
	#10 counter$count = 3660;
	#10 counter$count = 3661;
	#10 counter$count = 3662;
	#10 counter$count = 3663;
	#10 counter$count = 3664;
	#10 counter$count = 3665;
	#10 counter$count = 3666;
	#10 counter$count = 3667;
	#10 counter$count = 3668;
	#10 counter$count = 3669;
	#10 counter$count = 3670;
	#10 counter$count = 3671;
	#10 counter$count = 3672;
	#10 counter$count = 3673;
	#10 counter$count = 3674;
	#10 counter$count = 3675;
	#10 counter$count = 3676;
	#10 counter$count = 3677;
	#10 counter$count = 3678;
	#10 counter$count = 3679;
	#10 counter$count = 3680;
	#10 counter$count = 3681;
	#10 counter$count = 3682;
	#10 counter$count = 3683;
	#10 counter$count = 3684;
	#10 counter$count = 3685;
	#10 counter$count = 3686;
	#10 counter$count = 3687;
	#10 counter$count = 3688;
	#10 counter$count = 3689;
	#10 counter$count = 3690;
	#10 counter$count = 3691;
	#10 counter$count = 3692;
	#10 counter$count = 3693;
	#10 counter$count = 3694;
	#10 counter$count = 3695;
	#10 counter$count = 3696;
	#10 counter$count = 3697;
	#10 counter$count = 3698;
	#10 counter$count = 3699;
	#10 counter$count = 3700;
	#10 counter$count = 3701;
	#10 counter$count = 3702;
	#10 counter$count = 3703;
	#10 counter$count = 3704;
	#10 counter$count = 3705;
	#10 counter$count = 3706;
	#10 counter$count = 3707;
	#10 counter$count = 3708;
	#10 counter$count = 3709;
	#10 counter$count = 3710;
	#10 counter$count = 3711;
	#10 counter$count = 3712;
	#10 counter$count = 3713;
	#10 counter$count = 3714;
	#10 counter$count = 3715;
	#10 counter$count = 3716;
	#10 counter$count = 3717;
	#10 counter$count = 3718;
	#10 counter$count = 3719;
	#10 counter$count = 3720;
	#10 counter$count = 3721;
	#10 counter$count = 3722;
	#10 counter$count = 3723;
	#10 counter$count = 3724;
	#10 counter$count = 3725;
	#10 counter$count = 3726;
	#10 counter$count = 3727;
	#10 counter$count = 3728;
	#10 counter$count = 3729;
	#10 counter$count = 3730;
	#10 counter$count = 3731;
	#10 counter$count = 3732;
	#10 counter$count = 3733;
	#10 counter$count = 3734;
	#10 counter$count = 3735;
	#10 counter$count = 3736;
	#10 counter$count = 3737;
	#10 counter$count = 3738;
	#10 counter$count = 3739;
	#10 counter$count = 3740;
	#10 counter$count = 3741;
	#10 counter$count = 3742;
	#10 counter$count = 3743;
	#10 counter$count = 3744;
	#10 counter$count = 3745;
	#10 counter$count = 3746;
	#10 counter$count = 3747;
	#10 counter$count = 3748;
	#10 counter$count = 3749;
	#10 counter$count = 3750;
	#10 counter$count = 3751;
	#10 counter$count = 3752;
	#10 counter$count = 3753;
	#10 counter$count = 3754;
	#10 counter$count = 3755;
	#10 counter$count = 3756;
	#10 counter$count = 3757;
	#10 counter$count = 3758;
	#10 counter$count = 3759;
	#10 counter$count = 3760;
	#10 counter$count = 3761;
	#10 counter$count = 3762;
	#10 counter$count = 3763;
	#10 counter$count = 3764;
	#10 counter$count = 3765;
	#10 counter$count = 3766;
	#10 counter$count = 3767;
	#10 counter$count = 3768;
	#10 counter$count = 3769;
	#10 counter$count = 3770;
	#10 counter$count = 3771;
	#10 counter$count = 3772;
	#10 counter$count = 3773;
	#10 counter$count = 3774;
	#10 counter$count = 3775;
	#10 counter$count = 3776;
	#10 counter$count = 3777;
	#10 counter$count = 3778;
	#10 counter$count = 3779;
	#10 counter$count = 3780;
	#10 counter$count = 3781;
	#10 counter$count = 3782;
	#10 counter$count = 3783;
	#10 counter$count = 3784;
	#10 counter$count = 3785;
	#10 counter$count = 3786;
	#10 counter$count = 3787;
	#10 counter$count = 3788;
	#10 counter$count = 3789;
	#10 counter$count = 3790;
	#10 counter$count = 3791;
	#10 counter$count = 3792;
	#10 counter$count = 3793;
	#10 counter$count = 3794;
	#10 counter$count = 3795;
	#10 counter$count = 3796;
	#10 counter$count = 3797;
	#10 counter$count = 3798;
	#10 counter$count = 3799;
	#10 counter$count = 3800;
	#10 counter$count = 3801;
	#10 counter$count = 3802;
	#10 counter$count = 3803;
	#10 counter$count = 3804;
	#10 counter$count = 3805;
	#10 counter$count = 3806;
	#10 counter$count = 3807;
	#10 counter$count = 3808;
	#10 counter$count = 3809;
	#10 counter$count = 3810;
	#10 counter$count = 3811;
	#10 counter$count = 3812;
	#10 counter$count = 3813;
	#10 counter$count = 3814;
	#10 counter$count = 3815;
	#10 counter$count = 3816;
	#10 counter$count = 3817;
	#10 counter$count = 3818;
	#10 counter$count = 3819;
	#10 counter$count = 3820;
	#10 counter$count = 3821;
	#10 counter$count = 3822;
	#10 counter$count = 3823;
	#10 counter$count = 3824;
	#10 counter$count = 3825;
	#10 counter$count = 3826;
	#10 counter$count = 3827;
	#10 counter$count = 3828;
	#10 counter$count = 3829;
	#10 counter$count = 3830;
	#10 counter$count = 3831;
	#10 counter$count = 3832;
	#10 counter$count = 3833;
	#10 counter$count = 3834;
	#10 counter$count = 3835;
	#10 counter$count = 3836;
	#10 counter$count = 3837;
	#10 counter$count = 3838;
	#10 counter$count = 3839;
	#10 counter$count = 3840;
	#10 counter$count = 3841;
	#10 counter$count = 3842;
	#10 counter$count = 3843;
	#10 counter$count = 3844;
	#10 counter$count = 3845;
	#10 counter$count = 3846;
	#10 counter$count = 3847;
	#10 counter$count = 3848;
	#10 counter$count = 3849;
	#10 counter$count = 3850;
	#10 counter$count = 3851;
	#10 counter$count = 3852;
	#10 counter$count = 3853;
	#10 counter$count = 3854;
	#10 counter$count = 3855;
	#10 counter$count = 3856;
	#10 counter$count = 3857;
	#10 counter$count = 3858;
	#10 counter$count = 3859;
	#10 counter$count = 3860;
	#10 counter$count = 3861;
	#10 counter$count = 3862;
	#10 counter$count = 3863;
	#10 counter$count = 3864;
	#10 counter$count = 3865;
	#10 counter$count = 3866;
	#10 counter$count = 3867;
	#10 counter$count = 3868;
	#10 counter$count = 3869;
	#10 counter$count = 3870;
	#10 counter$count = 3871;
	#10 counter$count = 3872;
	#10 counter$count = 3873;
	#10 counter$count = 3874;
	#10 counter$count = 3875;
	#10 counter$count = 3876;
	#10 counter$count = 3877;
	#10 counter$count = 3878;
	#10 counter$count = 3879;
	#10 counter$count = 3880;
	#10 counter$count = 3881;
	#10 counter$count = 3882;
	#10 counter$count = 3883;
	#10 counter$count = 3884;
	#10 counter$count = 3885;
	#10 counter$count = 3886;
	#10 counter$count = 3887;
	#10 counter$count = 3888;
	#10 counter$count = 3889;
	#10 counter$count = 3890;
	#10 counter$count = 3891;
	#10 counter$count = 3892;
	#10 counter$count = 3893;
	#10 counter$count = 3894;
	#10 counter$count = 3895;
	#10 counter$count = 3896;
	#10 counter$count = 3897;
	#10 counter$count = 3898;
	#10 counter$count = 3899;
	#10 counter$count = 3900;
	#10 counter$count = 3901;
	#10 counter$count = 3902;
	#10 counter$count = 3903;
	#10 counter$count = 3904;
	#10 counter$count = 3905;
	#10 counter$count = 3906;
	#10 counter$count = 3907;
	#10 counter$count = 3908;
	#10 counter$count = 3909;
	#10 counter$count = 3910;
	#10 counter$count = 3911;
	#10 counter$count = 3912;
	#10 counter$count = 3913;
	#10 counter$count = 3914;
	#10 counter$count = 3915;
	#10 counter$count = 3916;
	#10 counter$count = 3917;
	#10 counter$count = 3918;
	#10 counter$count = 3919;
	#10 counter$count = 3920;
	#10 counter$count = 3921;
	#10 counter$count = 3922;
	#10 counter$count = 3923;
	#10 counter$count = 3924;
	#10 counter$count = 3925;
	#10 counter$count = 3926;
	#10 counter$count = 3927;
	#10 counter$count = 3928;
	#10 counter$count = 3929;
	#10 counter$count = 3930;
	#10 counter$count = 3931;
	#10 counter$count = 3932;
	#10 counter$count = 3933;
	#10 counter$count = 3934;
	#10 counter$count = 3935;
	#10 counter$count = 3936;
	#10 counter$count = 3937;
	#10 counter$count = 3938;
	#10 counter$count = 3939;
	#10 counter$count = 3940;
	#10 counter$count = 3941;
	#10 counter$count = 3942;
	#10 counter$count = 3943;
	#10 counter$count = 3944;
	#10 counter$count = 3945;
	#10 counter$count = 3946;
	#10 counter$count = 3947;
	#10 counter$count = 3948;
	#10 counter$count = 3949;
	#10 counter$count = 3950;
	#10 counter$count = 3951;
	#10 counter$count = 3952;
	#10 counter$count = 3953;
	#10 counter$count = 3954;
	#10 counter$count = 3955;
	#10 counter$count = 3956;
	#10 counter$count = 3957;
	#10 counter$count = 3958;
	#10 counter$count = 3959;
	#10 counter$count = 3960;
	#10 counter$count = 3961;
	#10 counter$count = 3962;
	#10 counter$count = 3963;
	#10 counter$count = 3964;
	#10 counter$count = 3965;
	#10 counter$count = 3966;
	#10 counter$count = 3967;
	#10 counter$count = 3968;
	#10 counter$count = 3969;
	#10 counter$count = 3970;
	#10 counter$count = 3971;
	#10 counter$count = 3972;
	#10 counter$count = 3973;
	#10 counter$count = 3974;
	#10 counter$count = 3975;
	#10 counter$count = 3976;
	#10 counter$count = 3977;
	#10 counter$count = 3978;
	#10 counter$count = 3979;
	#10 counter$count = 3980;
	#10 counter$count = 3981;
	#10 counter$count = 3982;
	#10 counter$count = 3983;
	#10 counter$count = 3984;
	#10 counter$count = 3985;
	#10 counter$count = 3986;
	#10 counter$count = 3987;
	#10 counter$count = 3988;
	#10 counter$count = 3989;
	#10 counter$count = 3990;
	#10 counter$count = 3991;
	#10 counter$count = 3992;
	#10 counter$count = 3993;
	#10 counter$count = 3994;
	#10 counter$count = 3995;
	#10 counter$count = 3996;
	#10 counter$count = 3997;
	#10 counter$count = 3998;
	#10 counter$count = 3999;
	#10 counter$count = 4000;
	#10 counter$count = 4001;
	#10 counter$count = 4002;
	#10 counter$count = 4003;
	#10 counter$count = 4004;
	#10 counter$count = 4005;
	#10 counter$count = 4006;
	#10 counter$count = 4007;
	#10 counter$count = 4008;
	#10 counter$count = 4009;
	#10 counter$count = 4010;
	#10 counter$count = 4011;
	#10 counter$count = 4012;
	#10 counter$count = 4013;
	#10 counter$count = 4014;
	#10 counter$count = 4015;
	#10 counter$count = 4016;
	#10 counter$count = 4017;
	#10 counter$count = 4018;
	#10 counter$count = 4019;
	#10 counter$count = 4020;
	#10 counter$count = 4021;
	#10 counter$count = 4022;
	#10 counter$count = 4023;
	#10 counter$count = 4024;
	#10 counter$count = 4025;
	#10 counter$count = 4026;
	#10 counter$count = 4027;
	#10 counter$count = 4028;
	#10 counter$count = 4029;
	#10 counter$count = 4030;
	#10 counter$count = 4031;
	#10 counter$count = 4032;
	#10 counter$count = 4033;
	#10 counter$count = 4034;
	#10 counter$count = 4035;
	#10 counter$count = 4036;
	#10 counter$count = 4037;
	#10 counter$count = 4038;
	#10 counter$count = 4039;
	#10 counter$count = 4040;
	#10 counter$count = 4041;
	#10 counter$count = 4042;
	#10 counter$count = 4043;
	#10 counter$count = 4044;
	#10 counter$count = 4045;
	#10 counter$count = 4046;
	#10 counter$count = 4047;
	#10 counter$count = 4048;
	#10 counter$count = 4049;
	#10 counter$count = 4050;
	#10 counter$count = 4051;
	#10 counter$count = 4052;
	#10 counter$count = 4053;
	#10 counter$count = 4054;
	#10 counter$count = 4055;
	#10 counter$count = 4056;
	#10 counter$count = 4057;
	#10 counter$count = 4058;
	#10 counter$count = 4059;
	#10 counter$count = 4060;
	#10 counter$count = 4061;
	#10 counter$count = 4062;
	#10 counter$count = 4063;
	#10 counter$count = 4064;
	#10 counter$count = 4065;
	#10 counter$count = 4066;
	#10 counter$count = 4067;
	#10 counter$count = 4068;
	#10 counter$count = 4069;
	#10 counter$count = 4070;
	#10 counter$count = 4071;
	#10 counter$count = 4072;
	#10 counter$count = 4073;
	#10 counter$count = 4074;
	#10 counter$count = 4075;
	#10 counter$count = 4076;
	#10 counter$count = 4077;
	#10 counter$count = 4078;
	#10 counter$count = 4079;
	#10 counter$count = 4080;
	#10 counter$count = 4081;
	#10 counter$count = 4082;
	#10 counter$count = 4083;
	#10 counter$count = 4084;
	#10 counter$count = 4085;
	#10 counter$count = 4086;
	#10 counter$count = 4087;
	#10 counter$count = 4088;
	#10 counter$count = 4089;
	#10 counter$count = 4090;
	#10 counter$count = 4091;
	#10 counter$count = 4092;
	#10 counter$count = 4093;
	#10 counter$count = 4094;
	#10 counter$count = 4095;
	#10 counter$count = 4096;
	#10 counter$count = 4097;
	#10 counter$count = 4098;
	#10 counter$count = 4099;
	#10 counter$count = 4100;
	#10 counter$count = 4101;
	#10 counter$count = 4102;
	#10 counter$count = 4103;
	#10 counter$count = 4104;
	#10 counter$count = 4105;
	#10 counter$count = 4106;
	#10 counter$count = 4107;
	#10 counter$count = 4108;
	#10 counter$count = 4109;
	#10 counter$count = 4110;
	#10 counter$count = 4111;
	#10 counter$count = 4112;
	#10 counter$count = 4113;
	#10 counter$count = 4114;
	#10 counter$count = 4115;
	#10 counter$count = 4116;
	#10 counter$count = 4117;
	#10 counter$count = 4118;
	#10 counter$count = 4119;
	#10 counter$count = 4120;
	#10 counter$count = 4121;
	#10 counter$count = 4122;
	#10 counter$count = 4123;
	#10 counter$count = 4124;
	#10 counter$count = 4125;
	#10 counter$count = 4126;
	#10 counter$count = 4127;
	#10 counter$count = 4128;
	#10 counter$count = 4129;
	#10 counter$count = 4130;
	#10 counter$count = 4131;
	#10 counter$count = 4132;
	#10 counter$count = 4133;
	#10 counter$count = 4134;
	#10 counter$count = 4135;
	#10 counter$count = 4136;
	#10 counter$count = 4137;
	#10 counter$count = 4138;
	#10 counter$count = 4139;
	#10 counter$count = 4140;
	#10 counter$count = 4141;
	#10 counter$count = 4142;
	#10 counter$count = 4143;
	#10 counter$count = 4144;
	#10 counter$count = 4145;
	#10 counter$count = 4146;
	#10 counter$count = 4147;
	#10 counter$count = 4148;
	#10 counter$count = 4149;
	#10 counter$count = 4150;
	#10 counter$count = 4151;
	#10 counter$count = 4152;
	#10 counter$count = 4153;
	#10 counter$count = 4154;
	#10 counter$count = 4155;
	#10 counter$count = 4156;
	#10 counter$count = 4157;
	#10 counter$count = 4158;
	#10 counter$count = 4159;
	#10 counter$count = 4160;
	#10 counter$count = 4161;
	#10 counter$count = 4162;
	#10 counter$count = 4163;
	#10 counter$count = 4164;
	#10 counter$count = 4165;
	#10 counter$count = 4166;
	#10 counter$count = 4167;
	#10 counter$count = 4168;
	#10 counter$count = 4169;
	#10 counter$count = 4170;
	#10 counter$count = 4171;
	#10 counter$count = 4172;
	#10 counter$count = 4173;
	#10 counter$count = 4174;
	#10 counter$count = 4175;
	#10 counter$count = 4176;
	#10 counter$count = 4177;
	#10 counter$count = 4178;
	#10 counter$count = 4179;
	#10 counter$count = 4180;
	#10 counter$count = 4181;
	#10 counter$count = 4182;
	#10 counter$count = 4183;
	#10 counter$count = 4184;
	#10 counter$count = 4185;
	#10 counter$count = 4186;
	#10 counter$count = 4187;
	#10 counter$count = 4188;
	#10 counter$count = 4189;
	#10 counter$count = 4190;
	#10 counter$count = 4191;
	#10 counter$count = 4192;
	#10 counter$count = 4193;
	#10 counter$count = 4194;
	#10 counter$count = 4195;
	#10 counter$count = 4196;
	#10 counter$count = 4197;
	#10 counter$count = 4198;
	#10 counter$count = 4199;
	#10 counter$count = 4200;
	#10 counter$count = 4201;
	#10 counter$count = 4202;
	#10 counter$count = 4203;
	#10 counter$count = 4204;
	#10 counter$count = 4205;
	#10 counter$count = 4206;
	#10 counter$count = 4207;
	#10 counter$count = 4208;
	#10 counter$count = 4209;
	#10 counter$count = 4210;
	#10 counter$count = 4211;
	#10 counter$count = 4212;
	#10 counter$count = 4213;
	#10 counter$count = 4214;
	#10 counter$count = 4215;
	#10 counter$count = 4216;
	#10 counter$count = 4217;
	#10 counter$count = 4218;
	#10 counter$count = 4219;
	#10 counter$count = 4220;
	#10 counter$count = 4221;
	#10 counter$count = 4222;
	#10 counter$count = 4223;
	#10 counter$count = 4224;
	#10 counter$count = 4225;
	#10 counter$count = 4226;
	#10 counter$count = 4227;
	#10 counter$count = 4228;
	#10 counter$count = 4229;
	#10 counter$count = 4230;
	#10 counter$count = 4231;
	#10 counter$count = 4232;
	#10 counter$count = 4233;
	#10 counter$count = 4234;
	#10 counter$count = 4235;
	#10 counter$count = 4236;
	#10 counter$count = 4237;
	#10 counter$count = 4238;
	#10 counter$count = 4239;
	#10 counter$count = 4240;
	#10 counter$count = 4241;
	#10 counter$count = 4242;
	#10 counter$count = 4243;
	#10 counter$count = 4244;
	#10 counter$count = 4245;
	#10 counter$count = 4246;
	#10 counter$count = 4247;
	#10 counter$count = 4248;
	#10 counter$count = 4249;
	#10 counter$count = 4250;
	#10 counter$count = 4251;
	#10 counter$count = 4252;
	#10 counter$count = 4253;
	#10 counter$count = 4254;
	#10 counter$count = 4255;
	#10 counter$count = 4256;
	#10 counter$count = 4257;
	#10 counter$count = 4258;
	#10 counter$count = 4259;
	#10 counter$count = 4260;
	#10 counter$count = 4261;
	#10 counter$count = 4262;
	#10 counter$count = 4263;
	#10 counter$count = 4264;
	#10 counter$count = 4265;
	#10 counter$count = 4266;
	#10 counter$count = 4267;
	#10 counter$count = 4268;
	#10 counter$count = 4269;
	#10 counter$count = 4270;
	#10 counter$count = 4271;
	#10 counter$count = 4272;
	#10 counter$count = 4273;
	#10 counter$count = 4274;
	#10 counter$count = 4275;
	#10 counter$count = 4276;
	#10 counter$count = 4277;
	#10 counter$count = 4278;
	#10 counter$count = 4279;
	#10 counter$count = 4280;
	#10 counter$count = 4281;
	#10 counter$count = 4282;
	#10 counter$count = 4283;
	#10 counter$count = 4284;
	#10 counter$count = 4285;
	#10 counter$count = 4286;
	#10 counter$count = 4287;
	#10 counter$count = 4288;
	#10 counter$count = 4289;
	#10 counter$count = 4290;
	#10 counter$count = 4291;
	#10 counter$count = 4292;
	#10 counter$count = 4293;
	#10 counter$count = 4294;
	#10 counter$count = 4295;
	#10 counter$count = 4296;
	#10 counter$count = 4297;
	#10 counter$count = 4298;
	#10 counter$count = 4299;
	#10 counter$count = 4300;
	#10 counter$count = 4301;
	#10 counter$count = 4302;
	#10 counter$count = 4303;
	#10 counter$count = 4304;
	#10 counter$count = 4305;
	#10 counter$count = 4306;
	#10 counter$count = 4307;
	#10 counter$count = 4308;
	#10 counter$count = 4309;
	#10 counter$count = 4310;
	#10 counter$count = 4311;
	#10 counter$count = 4312;
	#10 counter$count = 4313;
	#10 counter$count = 4314;
	#10 counter$count = 4315;
	#10 counter$count = 4316;
	#10 counter$count = 4317;
	#10 counter$count = 4318;
	#10 counter$count = 4319;
	#10 counter$count = 4320;
	#10 counter$count = 4321;
	#10 counter$count = 4322;
	#10 counter$count = 4323;
	#10 counter$count = 4324;
	#10 counter$count = 4325;
	#10 counter$count = 4326;
	#10 counter$count = 4327;
	#10 counter$count = 4328;
	#10 counter$count = 4329;
	#10 counter$count = 4330;
	#10 counter$count = 4331;
	#10 counter$count = 4332;
	#10 counter$count = 4333;
	#10 counter$count = 4334;
	#10 counter$count = 4335;
	#10 counter$count = 4336;
	#10 counter$count = 4337;
	#10 counter$count = 4338;
	#10 counter$count = 4339;
	#10 counter$count = 4340;
	#10 counter$count = 4341;
	#10 counter$count = 4342;
	#10 counter$count = 4343;
	#10 counter$count = 4344;
	#10 counter$count = 4345;
	#10 counter$count = 4346;
	#10 counter$count = 4347;
	#10 counter$count = 4348;
	#10 counter$count = 4349;
	#10 counter$count = 4350;
	#10 counter$count = 4351;
	#10 counter$count = 4352;
	#10 counter$count = 4353;
	#10 counter$count = 4354;
	#10 counter$count = 4355;
	#10 counter$count = 4356;
	#10 counter$count = 4357;
	#10 counter$count = 4358;
	#10 counter$count = 4359;
	#10 counter$count = 4360;
	#10 counter$count = 4361;
	#10 counter$count = 4362;
	#10 counter$count = 4363;
	#10 counter$count = 4364;
	#10 counter$count = 4365;
	#10 counter$count = 4366;
	#10 counter$count = 4367;
	#10 counter$count = 4368;
	#10 counter$count = 4369;
	#10 counter$count = 4370;
	#10 counter$count = 4371;
	#10 counter$count = 4372;
	#10 counter$count = 4373;
	#10 counter$count = 4374;
	#10 counter$count = 4375;
	#10 counter$count = 4376;
	#10 counter$count = 4377;
	#10 counter$count = 4378;
	#10 counter$count = 4379;
	#10 counter$count = 4380;
	#10 counter$count = 4381;
	#10 counter$count = 4382;
	#10 counter$count = 4383;
	#10 counter$count = 4384;
	#10 counter$count = 4385;
	#10 counter$count = 4386;
	#10 counter$count = 4387;
	#10 counter$count = 4388;
	#10 counter$count = 4389;
	#10 counter$count = 4390;
	#10 counter$count = 4391;
	#10 counter$count = 4392;
	#10 counter$count = 4393;
	#10 counter$count = 4394;
	#10 counter$count = 4395;
	#10 counter$count = 4396;
	#10 counter$count = 4397;
	#10 counter$count = 4398;
	#10 counter$count = 4399;
	#10 counter$count = 4400;
	#10 counter$count = 4401;
	#10 counter$count = 4402;
	#10 counter$count = 4403;
	#10 counter$count = 4404;
	#10 counter$count = 4405;
	#10 counter$count = 4406;
	#10 counter$count = 4407;
	#10 counter$count = 4408;
	#10 counter$count = 4409;
	#10 counter$count = 4410;
	#10 counter$count = 4411;
	#10 counter$count = 4412;
	#10 counter$count = 4413;
	#10 counter$count = 4414;
	#10 counter$count = 4415;
	#10 counter$count = 4416;
	#10 counter$count = 4417;
	#10 counter$count = 4418;
	#10 counter$count = 4419;
	#10 counter$count = 4420;
	#10 counter$count = 4421;
	#10 counter$count = 4422;
	#10 counter$count = 4423;
	#10 counter$count = 4424;
	#10 counter$count = 4425;
	#10 counter$count = 4426;
	#10 counter$count = 4427;
	#10 counter$count = 4428;
	#10 counter$count = 4429;
	#10 counter$count = 4430;
	#10 counter$count = 4431;
	#10 counter$count = 4432;
	#10 counter$count = 4433;
	#10 counter$count = 4434;
	#10 counter$count = 4435;
	#10 counter$count = 4436;
	#10 counter$count = 4437;
	#10 counter$count = 4438;
	#10 counter$count = 4439;
	#10 counter$count = 4440;
	#10 counter$count = 4441;
	#10 counter$count = 4442;
	#10 counter$count = 4443;
	#10 counter$count = 4444;
	#10 counter$count = 4445;
	#10 counter$count = 4446;
	#10 counter$count = 4447;
	#10 counter$count = 4448;
	#10 counter$count = 4449;
	#10 counter$count = 4450;
	#10 counter$count = 4451;
	#10 counter$count = 4452;
	#10 counter$count = 4453;
	#10 counter$count = 4454;
	#10 counter$count = 4455;
	#10 counter$count = 4456;
	#10 counter$count = 4457;
	#10 counter$count = 4458;
	#10 counter$count = 4459;
	#10 counter$count = 4460;
	#10 counter$count = 4461;
	#10 counter$count = 4462;
	#10 counter$count = 4463;
	#10 counter$count = 4464;
	#10 counter$count = 4465;
	#10 counter$count = 4466;
	#10 counter$count = 4467;
	#10 counter$count = 4468;
	#10 counter$count = 4469;
	#10 counter$count = 4470;
	#10 counter$count = 4471;
	#10 counter$count = 4472;
	#10 counter$count = 4473;
	#10 counter$count = 4474;
	#10 counter$count = 4475;
	#10 counter$count = 4476;
	#10 counter$count = 4477;
	#10 counter$count = 4478;
	#10 counter$count = 4479;
	#10 counter$count = 4480;
	#10 counter$count = 4481;
	#10 counter$count = 4482;
	#10 counter$count = 4483;
	#10 counter$count = 4484;
	#10 counter$count = 4485;
	#10 counter$count = 4486;
	#10 counter$count = 4487;
	#10 counter$count = 4488;
	#10 counter$count = 4489;
	#10 counter$count = 4490;
	#10 counter$count = 4491;
	#10 counter$count = 4492;
	#10 counter$count = 4493;
	#10 counter$count = 4494;
	#10 counter$count = 4495;
	#10 counter$count = 4496;
	#10 counter$count = 4497;
	#10 counter$count = 4498;
	#10 counter$count = 4499;
	#10 counter$count = 4500;
	#10 counter$count = 4501;
	#10 counter$count = 4502;
	#10 counter$count = 4503;
	#10 counter$count = 4504;
	#10 counter$count = 4505;
	#10 counter$count = 4506;
	#10 counter$count = 4507;
	#10 counter$count = 4508;
	#10 counter$count = 4509;
	#10 counter$count = 4510;
	#10 counter$count = 4511;
	#10 counter$count = 4512;
	#10 counter$count = 4513;
	#10 counter$count = 4514;
	#10 counter$count = 4515;
	#10 counter$count = 4516;
	#10 counter$count = 4517;
	#10 counter$count = 4518;
	#10 counter$count = 4519;
	#10 counter$count = 4520;
	#10 counter$count = 4521;
	#10 counter$count = 4522;
	#10 counter$count = 4523;
	#10 counter$count = 4524;
	#10 counter$count = 4525;
	#10 counter$count = 4526;
	#10 counter$count = 4527;
	#10 counter$count = 4528;
	#10 counter$count = 4529;
	#10 counter$count = 4530;
	#10 counter$count = 4531;
	#10 counter$count = 4532;
	#10 counter$count = 4533;
	#10 counter$count = 4534;
	#10 counter$count = 4535;
	#10 counter$count = 4536;
	#10 counter$count = 4537;
	#10 counter$count = 4538;
	#10 counter$count = 4539;
	#10 counter$count = 4540;
	#10 counter$count = 4541;
	#10 counter$count = 4542;
	#10 counter$count = 4543;
	#10 counter$count = 4544;
	#10 counter$count = 4545;
	#10 counter$count = 4546;
	#10 counter$count = 4547;
	#10 counter$count = 4548;
	#10 counter$count = 4549;
	#10 counter$count = 4550;
	#10 counter$count = 4551;
	#10 counter$count = 4552;
	#10 counter$count = 4553;
	#10 counter$count = 4554;
	#10 counter$count = 4555;
	#10 counter$count = 4556;
	#10 counter$count = 4557;
	#10 counter$count = 4558;
	#10 counter$count = 4559;
	#10 counter$count = 4560;
	#10 counter$count = 4561;
	#10 counter$count = 4562;
	#10 counter$count = 4563;
	#10 counter$count = 4564;
	#10 counter$count = 4565;
	#10 counter$count = 4566;
	#10 counter$count = 4567;
	#10 counter$count = 4568;
	#10 counter$count = 4569;
	#10 counter$count = 4570;
	#10 counter$count = 4571;
	#10 counter$count = 4572;
	#10 counter$count = 4573;
	#10 counter$count = 4574;
	#10 counter$count = 4575;
	#10 counter$count = 4576;
	#10 counter$count = 4577;
	#10 counter$count = 4578;
	#10 counter$count = 4579;
	#10 counter$count = 4580;
	#10 counter$count = 4581;
	#10 counter$count = 4582;
	#10 counter$count = 4583;
	#10 counter$count = 4584;
	#10 counter$count = 4585;
	#10 counter$count = 4586;
	#10 counter$count = 4587;
	#10 counter$count = 4588;
	#10 counter$count = 4589;
	#10 counter$count = 4590;
	#10 counter$count = 4591;
	#10 counter$count = 4592;
	#10 counter$count = 4593;
	#10 counter$count = 4594;
	#10 counter$count = 4595;
	#10 counter$count = 4596;
	#10 counter$count = 4597;
	#10 counter$count = 4598;
	#10 counter$count = 4599;
	#10 counter$count = 4600;
	#10 counter$count = 4601;
	#10 counter$count = 4602;
	#10 counter$count = 4603;
	#10 counter$count = 4604;
	#10 counter$count = 4605;
	#10 counter$count = 4606;
	#10 counter$count = 4607;
	#10 counter$count = 4608;
	#10 counter$count = 4609;
	#10 counter$count = 4610;
	#10 counter$count = 4611;
	#10 counter$count = 4612;
	#10 counter$count = 4613;
	#10 counter$count = 4614;
	#10 counter$count = 4615;
	#10 counter$count = 4616;
	#10 counter$count = 4617;
	#10 counter$count = 4618;
	#10 counter$count = 4619;
	#10 counter$count = 4620;
	#10 counter$count = 4621;
	#10 counter$count = 4622;
	#10 counter$count = 4623;
	#10 counter$count = 4624;
	#10 counter$count = 4625;
	#10 counter$count = 4626;
	#10 counter$count = 4627;
	#10 counter$count = 4628;
	#10 counter$count = 4629;
	#10 counter$count = 4630;
	#10 counter$count = 4631;
	#10 counter$count = 4632;
	#10 counter$count = 4633;
	#10 counter$count = 4634;
	#10 counter$count = 4635;
	#10 counter$count = 4636;
	#10 counter$count = 4637;
	#10 counter$count = 4638;
	#10 counter$count = 4639;
	#10 counter$count = 4640;
	#10 counter$count = 4641;
	#10 counter$count = 4642;
	#10 counter$count = 4643;
	#10 counter$count = 4644;
	#10 counter$count = 4645;
	#10 counter$count = 4646;
	#10 counter$count = 4647;
	#10 counter$count = 4648;
	#10 counter$count = 4649;
	#10 counter$count = 4650;
	#10 counter$count = 4651;
	#10 counter$count = 4652;
	#10 counter$count = 4653;
	#10 counter$count = 4654;
	#10 counter$count = 4655;
	#10 counter$count = 4656;
	#10 counter$count = 4657;
	#10 counter$count = 4658;
	#10 counter$count = 4659;
	#10 counter$count = 4660;
	#10 counter$count = 4661;
	#10 counter$count = 4662;
	#10 counter$count = 4663;
	#10 counter$count = 4664;
	#10 counter$count = 4665;
	#10 counter$count = 4666;
	#10 counter$count = 4667;
	#10 counter$count = 4668;
	#10 counter$count = 4669;
	#10 counter$count = 4670;
	#10 counter$count = 4671;
	#10 counter$count = 4672;
	#10 counter$count = 4673;
	#10 counter$count = 4674;
	#10 counter$count = 4675;
	#10 counter$count = 4676;
	#10 counter$count = 4677;
	#10 counter$count = 4678;
	#10 counter$count = 4679;
	#10 counter$count = 4680;
	#10 counter$count = 4681;
	#10 counter$count = 4682;
	#10 counter$count = 4683;
	#10 counter$count = 4684;
	#10 counter$count = 4685;
	#10 counter$count = 4686;
	#10 counter$count = 4687;
	#10 counter$count = 4688;
	#10 counter$count = 4689;
	#10 counter$count = 4690;
	#10 counter$count = 4691;
	#10 counter$count = 4692;
	#10 counter$count = 4693;
	#10 counter$count = 4694;
	#10 counter$count = 4695;
	#10 counter$count = 4696;
	#10 counter$count = 4697;
	#10 counter$count = 4698;
	#10 counter$count = 4699;
	#10 counter$count = 4700;
	#10 counter$count = 4701;
	#10 counter$count = 4702;
	#10 counter$count = 4703;
	#10 counter$count = 4704;
	#10 counter$count = 4705;
	#10 counter$count = 4706;
	#10 counter$count = 4707;
	#10 counter$count = 4708;
	#10 counter$count = 4709;
	#10 counter$count = 4710;
	#10 counter$count = 4711;
	#10 counter$count = 4712;
	#10 counter$count = 4713;
	#10 counter$count = 4714;
	#10 counter$count = 4715;
	#10 counter$count = 4716;
	#10 counter$count = 4717;
	#10 counter$count = 4718;
	#10 counter$count = 4719;
	#10 counter$count = 4720;
	#10 counter$count = 4721;
	#10 counter$count = 4722;
	#10 counter$count = 4723;
	#10 counter$count = 4724;
	#10 counter$count = 4725;
	#10 counter$count = 4726;
	#10 counter$count = 4727;
	#10 counter$count = 4728;
	#10 counter$count = 4729;
	#10 counter$count = 4730;
	#10 counter$count = 4731;
	#10 counter$count = 4732;
	#10 counter$count = 4733;
	#10 counter$count = 4734;
	#10 counter$count = 4735;
	#10 counter$count = 4736;
	#10 counter$count = 4737;
	#10 counter$count = 4738;
	#10 counter$count = 4739;
	#10 counter$count = 4740;
	#10 counter$count = 4741;
	#10 counter$count = 4742;
	#10 counter$count = 4743;
	#10 counter$count = 4744;
	#10 counter$count = 4745;
	#10 counter$count = 4746;
	#10 counter$count = 4747;
	#10 counter$count = 4748;
	#10 counter$count = 4749;
	#10 counter$count = 4750;
	#10 counter$count = 4751;
	#10 counter$count = 4752;
	#10 counter$count = 4753;
	#10 counter$count = 4754;
	#10 counter$count = 4755;
	#10 counter$count = 4756;
	#10 counter$count = 4757;
	#10 counter$count = 4758;
	#10 counter$count = 4759;
	#10 counter$count = 4760;
	#10 counter$count = 4761;
	#10 counter$count = 4762;
	#10 counter$count = 4763;
	#10 counter$count = 4764;
	#10 counter$count = 4765;
	#10 counter$count = 4766;
	#10 counter$count = 4767;
	#10 counter$count = 4768;
	#10 counter$count = 4769;
	#10 counter$count = 4770;
	#10 counter$count = 4771;
	#10 counter$count = 4772;
	#10 counter$count = 4773;
	#10 counter$count = 4774;
	#10 counter$count = 4775;
	#10 counter$count = 4776;
	#10 counter$count = 4777;
	#10 counter$count = 4778;
	#10 counter$count = 4779;
	#10 counter$count = 4780;
	#10 counter$count = 4781;
	#10 counter$count = 4782;
	#10 counter$count = 4783;
	#10 counter$count = 4784;
	#10 counter$count = 4785;
	#10 counter$count = 4786;
	#10 counter$count = 4787;
	#10 counter$count = 4788;
	#10 counter$count = 4789;
	#10 counter$count = 4790;
	#10 counter$count = 4791;
	#10 counter$count = 4792;
	#10 counter$count = 4793;
	#10 counter$count = 4794;
	#10 counter$count = 4795;
	#10 counter$count = 4796;
	#10 counter$count = 4797;
	#10 counter$count = 4798;
	#10 counter$count = 4799;
	#10 counter$count = 4800;
	#10 counter$count = 4801;
	#10 counter$count = 4802;
	#10 counter$count = 4803;
	#10 counter$count = 4804;
	#10 counter$count = 4805;
	#10 counter$count = 4806;
	#10 counter$count = 4807;
	#10 counter$count = 4808;
	#10 counter$count = 4809;
	#10 counter$count = 4810;
	#10 counter$count = 4811;
	#10 counter$count = 4812;
	#10 counter$count = 4813;
	#10 counter$count = 4814;
	#10 counter$count = 4815;
	#10 counter$count = 4816;
	#10 counter$count = 4817;
	#10 counter$count = 4818;
	#10 counter$count = 4819;
	#10 counter$count = 4820;
	#10 counter$count = 4821;
	#10 counter$count = 4822;
	#10 counter$count = 4823;
	#10 counter$count = 4824;
	#10 counter$count = 4825;
	#10 counter$count = 4826;
	#10 counter$count = 4827;
	#10 counter$count = 4828;
	#10 counter$count = 4829;
	#10 counter$count = 4830;
	#10 counter$count = 4831;
	#10 counter$count = 4832;
	#10 counter$count = 4833;
	#10 counter$count = 4834;
	#10 counter$count = 4835;
	#10 counter$count = 4836;
	#10 counter$count = 4837;
	#10 counter$count = 4838;
	#10 counter$count = 4839;
	#10 counter$count = 4840;
	#10 counter$count = 4841;
	#10 counter$count = 4842;
	#10 counter$count = 4843;
	#10 counter$count = 4844;
	#10 counter$count = 4845;
	#10 counter$count = 4846;
	#10 counter$count = 4847;
	#10 counter$count = 4848;
	#10 counter$count = 4849;
	#10 counter$count = 4850;
	#10 counter$count = 4851;
	#10 counter$count = 4852;
	#10 counter$count = 4853;
	#10 counter$count = 4854;
	#10 counter$count = 4855;
	#10 counter$count = 4856;
	#10 counter$count = 4857;
	#10 counter$count = 4858;
	#10 counter$count = 4859;
	#10 counter$count = 4860;
	#10 counter$count = 4861;
	#10 counter$count = 4862;
	#10 counter$count = 4863;
	#10 counter$count = 4864;
	#10 counter$count = 4865;
	#10 counter$count = 4866;
	#10 counter$count = 4867;
	#10 counter$count = 4868;
	#10 counter$count = 4869;
	#10 counter$count = 4870;
	#10 counter$count = 4871;
	#10 counter$count = 4872;
	#10 counter$count = 4873;
	#10 counter$count = 4874;
	#10 counter$count = 4875;
	#10 counter$count = 4876;
	#10 counter$count = 4877;
	#10 counter$count = 4878;
	#10 counter$count = 4879;
	#10 counter$count = 4880;
	#10 counter$count = 4881;
	#10 counter$count = 4882;
	#10 counter$count = 4883;
	#10 counter$count = 4884;
	#10 counter$count = 4885;
	#10 counter$count = 4886;
	#10 counter$count = 4887;
	#10 counter$count = 4888;
	#10 counter$count = 4889;
	#10 counter$count = 4890;
	#10 counter$count = 4891;
	#10 counter$count = 4892;
	#10 counter$count = 4893;
	#10 counter$count = 4894;
	#10 counter$count = 4895;
	#10 counter$count = 4896;
	#10 counter$count = 4897;
	#10 counter$count = 4898;
	#10 counter$count = 4899;
	#10 counter$count = 4900;
	#10 counter$count = 4901;
	#10 counter$count = 4902;
	#10 counter$count = 4903;
	#10 counter$count = 4904;
	#10 counter$count = 4905;
	#10 counter$count = 4906;
	#10 counter$count = 4907;
	#10 counter$count = 4908;
	#10 counter$count = 4909;
	#10 counter$count = 4910;
	#10 counter$count = 4911;
	#10 counter$count = 4912;
	#10 counter$count = 4913;
	#10 counter$count = 4914;
	#10 counter$count = 4915;
	#10 counter$count = 4916;
	#10 counter$count = 4917;
	#10 counter$count = 4918;
	#10 counter$count = 4919;
	#10 counter$count = 4920;
	#10 counter$count = 4921;
	#10 counter$count = 4922;
	#10 counter$count = 4923;
	#10 counter$count = 4924;
	#10 counter$count = 4925;
	#10 counter$count = 4926;
	#10 counter$count = 4927;
	#10 counter$count = 4928;
	#10 counter$count = 4929;
	#10 counter$count = 4930;
	#10 counter$count = 4931;
	#10 counter$count = 4932;
	#10 counter$count = 4933;
	#10 counter$count = 4934;
	#10 counter$count = 4935;
	#10 counter$count = 4936;
	#10 counter$count = 4937;
	#10 counter$count = 4938;
	#10 counter$count = 4939;
	#10 counter$count = 4940;
	#10 counter$count = 4941;
	#10 counter$count = 4942;
	#10 counter$count = 4943;
	#10 counter$count = 4944;
	#10 counter$count = 4945;
	#10 counter$count = 4946;
	#10 counter$count = 4947;
	#10 counter$count = 4948;
	#10 counter$count = 4949;
	#10 counter$count = 4950;
	#10 counter$count = 4951;
	#10 counter$count = 4952;
	#10 counter$count = 4953;
	#10 counter$count = 4954;
	#10 counter$count = 4955;
	#10 counter$count = 4956;
	#10 counter$count = 4957;
	#10 counter$count = 4958;
	#10 counter$count = 4959;
	#10 counter$count = 4960;
	#10 counter$count = 4961;
	#10 counter$count = 4962;
	#10 counter$count = 4963;
	#10 counter$count = 4964;
	#10 counter$count = 4965;
	#10 counter$count = 4966;
	#10 counter$count = 4967;
	#10 counter$count = 4968;
	#10 counter$count = 4969;
	#10 counter$count = 4970;
	#10 counter$count = 4971;
	#10 counter$count = 4972;
	#10 counter$count = 4973;
	#10 counter$count = 4974;
	#10 counter$count = 4975;
	#10 counter$count = 4976;
	#10 counter$count = 4977;
	#10 counter$count = 4978;
	#10 counter$count = 4979;
	#10 counter$count = 4980;
	#10 counter$count = 4981;
	#10 counter$count = 4982;
	#10 counter$count = 4983;
	#10 counter$count = 4984;
	#10 counter$count = 4985;
	#10 counter$count = 4986;
	#10 counter$count = 4987;
	#10 counter$count = 4988;
	#10 counter$count = 4989;
	#10 counter$count = 4990;
	#10 counter$count = 4991;
	#10 counter$count = 4992;
	#10 counter$count = 4993;
	#10 counter$count = 4994;
	#10 counter$count = 4995;
	#10 counter$count = 4996;
	#10 counter$count = 4997;
	#10 counter$count = 4998;
	#10 counter$count = 4999;
	#10 counter$count = 5000;
	#10 counter$count = 5001;
	#10 counter$count = 5002;
	#10 counter$count = 5003;
	#10 counter$count = 5004;
	#10 counter$count = 5005;
	#10 counter$count = 5006;
	#10 counter$count = 5007;
	#10 counter$count = 5008;
	#10 counter$count = 5009;
	#10 counter$count = 5010;
	#10 counter$count = 5011;
	#10 counter$count = 5012;
	#10 counter$count = 5013;
	#10 counter$count = 5014;
	#10 counter$count = 5015;
	#10 counter$count = 5016;
	#10 counter$count = 5017;
	#10 counter$count = 5018;
	#10 counter$count = 5019;
	#10 counter$count = 5020;
	#10 counter$count = 5021;
	#10 counter$count = 5022;
	#10 counter$count = 5023;
	#10 counter$count = 5024;
	#10 counter$count = 5025;
	#10 counter$count = 5026;
	#10 counter$count = 5027;
	#10 counter$count = 5028;
	#10 counter$count = 5029;
	#10 counter$count = 5030;
	#10 counter$count = 5031;
	#10 counter$count = 5032;
	#10 counter$count = 5033;
	#10 counter$count = 5034;
	#10 counter$count = 5035;
	#10 counter$count = 5036;
	#10 counter$count = 5037;
	#10 counter$count = 5038;
	#10 counter$count = 5039;
	#10 counter$count = 5040;
	#10 counter$count = 5041;
	#10 counter$count = 5042;
	#10 counter$count = 5043;
	#10 counter$count = 5044;
	#10 counter$count = 5045;
	#10 counter$count = 5046;
	#10 counter$count = 5047;
	#10 counter$count = 5048;
	#10 counter$count = 5049;
	#10 counter$count = 5050;
	#10 counter$count = 5051;
	#10 counter$count = 5052;
	#10 counter$count = 5053;
	#10 counter$count = 5054;
	#10 counter$count = 5055;
	#10 counter$count = 5056;
	#10 counter$count = 5057;
	#10 counter$count = 5058;
	#10 counter$count = 5059;
	#10 counter$count = 5060;
	#10 counter$count = 5061;
	#10 counter$count = 5062;
	#10 counter$count = 5063;
	#10 counter$count = 5064;
	#10 counter$count = 5065;
	#10 counter$count = 5066;
	#10 counter$count = 5067;
	#10 counter$count = 5068;
	#10 counter$count = 5069;
	#10 counter$count = 5070;
	#10 counter$count = 5071;
	#10 counter$count = 5072;
	#10 counter$count = 5073;
	#10 counter$count = 5074;
	#10 counter$count = 5075;
	#10 counter$count = 5076;
	#10 counter$count = 5077;
	#10 counter$count = 5078;
	#10 counter$count = 5079;
	#10 counter$count = 5080;
	#10 counter$count = 5081;
	#10 counter$count = 5082;
	#10 counter$count = 5083;
	#10 counter$count = 5084;
	#10 counter$count = 5085;
	#10 counter$count = 5086;
	#10 counter$count = 5087;
	#10 counter$count = 5088;
	#10 counter$count = 5089;
	#10 counter$count = 5090;
	#10 counter$count = 5091;
	#10 counter$count = 5092;
	#10 counter$count = 5093;
	#10 counter$count = 5094;
	#10 counter$count = 5095;
	#10 counter$count = 5096;
	#10 counter$count = 5097;
	#10 counter$count = 5098;
	#10 counter$count = 5099;
	#10 counter$count = 5100;
	#10 counter$count = 5101;
	#10 counter$count = 5102;
	#10 counter$count = 5103;
	#10 counter$count = 5104;
	#10 counter$count = 5105;
	#10 counter$count = 5106;
	#10 counter$count = 5107;
	#10 counter$count = 5108;
	#10 counter$count = 5109;
	#10 counter$count = 5110;
	#10 counter$count = 5111;
	#10 counter$count = 5112;
	#10 counter$count = 5113;
	#10 counter$count = 5114;
	#10 counter$count = 5115;
	#10 counter$count = 5116;
	#10 counter$count = 5117;
	#10 counter$count = 5118;
	#10 counter$count = 5119;
	#10 counter$count = 5120;
	#10 counter$count = 5121;
	#10 counter$count = 5122;
	#10 counter$count = 5123;
	#10 counter$count = 5124;
	#10 counter$count = 5125;
	#10 counter$count = 5126;
	#10 counter$count = 5127;
	#10 counter$count = 5128;
	#10 counter$count = 5129;
	#10 counter$count = 5130;
	#10 counter$count = 5131;
	#10 counter$count = 5132;
	#10 counter$count = 5133;
	#10 counter$count = 5134;
	#10 counter$count = 5135;
	#10 counter$count = 5136;
	#10 counter$count = 5137;
	#10 counter$count = 5138;
	#10 counter$count = 5139;
	#10 counter$count = 5140;
	#10 counter$count = 5141;
	#10 counter$count = 5142;
	#10 counter$count = 5143;
	#10 counter$count = 5144;
	#10 counter$count = 5145;
	#10 counter$count = 5146;
	#10 counter$count = 5147;
	#10 counter$count = 5148;
	#10 counter$count = 5149;
	#10 counter$count = 5150;
	#10 counter$count = 5151;
	#10 counter$count = 5152;
	#10 counter$count = 5153;
	#10 counter$count = 5154;
	#10 counter$count = 5155;
	#10 counter$count = 5156;
	#10 counter$count = 5157;
	#10 counter$count = 5158;
	#10 counter$count = 5159;
	#10 counter$count = 5160;
	#10 counter$count = 5161;
	#10 counter$count = 5162;
	#10 counter$count = 5163;
	#10 counter$count = 5164;
	#10 counter$count = 5165;
	#10 counter$count = 5166;
	#10 counter$count = 5167;
	#10 counter$count = 5168;
	#10 counter$count = 5169;
	#10 counter$count = 5170;
	#10 counter$count = 5171;
	#10 counter$count = 5172;
	#10 counter$count = 5173;
	#10 counter$count = 5174;
	#10 counter$count = 5175;
	#10 counter$count = 5176;
	#10 counter$count = 5177;
	#10 counter$count = 5178;
	#10 counter$count = 5179;
	#10 counter$count = 5180;
	#10 counter$count = 5181;
	#10 counter$count = 5182;
	#10 counter$count = 5183;
	#10 counter$count = 5184;
	#10 counter$count = 5185;
	#10 counter$count = 5186;
	#10 counter$count = 5187;
	#10 counter$count = 5188;
	#10 counter$count = 5189;
	#10 counter$count = 5190;
	#10 counter$count = 5191;
	#10 counter$count = 5192;
	#10 counter$count = 5193;
	#10 counter$count = 5194;
	#10 counter$count = 5195;
	#10 counter$count = 5196;
	#10 counter$count = 5197;
	#10 counter$count = 5198;
	#10 counter$count = 5199;
	#10 counter$count = 5200;
	#10 counter$count = 5201;
	#10 counter$count = 5202;
	#10 counter$count = 5203;
	#10 counter$count = 5204;
	#10 counter$count = 5205;
	#10 counter$count = 5206;
	#10 counter$count = 5207;
	#10 counter$count = 5208;
	#10 counter$count = 5209;
	#10 counter$count = 5210;
	#10 counter$count = 5211;
	#10 counter$count = 5212;
	#10 counter$count = 5213;
	#10 counter$count = 5214;
	#10 counter$count = 5215;
	#10 counter$count = 5216;
	#10 counter$count = 5217;
	#10 counter$count = 5218;
	#10 counter$count = 5219;
	#10 counter$count = 5220;
	#10 counter$count = 5221;
	#10 counter$count = 5222;
	#10 counter$count = 5223;
	#10 counter$count = 5224;
	#10 counter$count = 5225;
	#10 counter$count = 5226;
	#10 counter$count = 5227;
	#10 counter$count = 5228;
	#10 counter$count = 5229;
	#10 counter$count = 5230;
	#10 counter$count = 5231;
	#10 counter$count = 5232;
	#10 counter$count = 5233;
	#10 counter$count = 5234;
	#10 counter$count = 5235;
	#10 counter$count = 5236;
	#10 counter$count = 5237;
	#10 counter$count = 5238;
	#10 counter$count = 5239;
	#10 counter$count = 5240;
	#10 counter$count = 5241;
	#10 counter$count = 5242;
	#10 counter$count = 5243;
	#10 counter$count = 5244;
	#10 counter$count = 5245;
	#10 counter$count = 5246;
	#10 counter$count = 5247;
	#10 counter$count = 5248;
	#10 counter$count = 5249;
	#10 counter$count = 5250;
	#10 counter$count = 5251;
	#10 counter$count = 5252;
	#10 counter$count = 5253;
	#10 counter$count = 5254;
	#10 counter$count = 5255;
	#10 counter$count = 5256;
	#10 counter$count = 5257;
	#10 counter$count = 5258;
	#10 counter$count = 5259;
	#10 counter$count = 5260;
	#10 counter$count = 5261;
	#10 counter$count = 5262;
	#10 counter$count = 5263;
	#10 counter$count = 5264;
	#10 counter$count = 5265;
	#10 counter$count = 5266;
	#10 counter$count = 5267;
	#10 counter$count = 5268;
	#10 counter$count = 5269;
	#10 counter$count = 5270;
	#10 counter$count = 5271;
	#10 counter$count = 5272;
	#10 counter$count = 5273;
	#10 counter$count = 5274;
	#10 counter$count = 5275;
	#10 counter$count = 5276;
	#10 counter$count = 5277;
	#10 counter$count = 5278;
	#10 counter$count = 5279;
	#10 counter$count = 5280;
	#10 counter$count = 5281;
	#10 counter$count = 5282;
	#10 counter$count = 5283;
	#10 counter$count = 5284;
	#10 counter$count = 5285;
	#10 counter$count = 5286;
	#10 counter$count = 5287;
	#10 counter$count = 5288;
	#10 counter$count = 5289;
	#10 counter$count = 5290;
	#10 counter$count = 5291;
	#10 counter$count = 5292;
	#10 counter$count = 5293;
	#10 counter$count = 5294;
	#10 counter$count = 5295;
	#10 counter$count = 5296;
	#10 counter$count = 5297;
	#10 counter$count = 5298;
	#10 counter$count = 5299;
	#10 counter$count = 5300;
	#10 counter$count = 5301;
	#10 counter$count = 5302;
	#10 counter$count = 5303;
	#10 counter$count = 5304;
	#10 counter$count = 5305;
	#10 counter$count = 5306;
	#10 counter$count = 5307;
	#10 counter$count = 5308;
	#10 counter$count = 5309;
	#10 counter$count = 5310;
	#10 counter$count = 5311;
	#10 counter$count = 5312;
	#10 counter$count = 5313;
	#10 counter$count = 5314;
	#10 counter$count = 5315;
	#10 counter$count = 5316;
	#10 counter$count = 5317;
	#10 counter$count = 5318;
	#10 counter$count = 5319;
	#10 counter$count = 5320;
	#10 counter$count = 5321;
	#10 counter$count = 5322;
	#10 counter$count = 5323;
	#10 counter$count = 5324;
	#10 counter$count = 5325;
	#10 counter$count = 5326;
	#10 counter$count = 5327;
	#10 counter$count = 5328;
	#10 counter$count = 5329;
	#10 counter$count = 5330;
	#10 counter$count = 5331;
	#10 counter$count = 5332;
	#10 counter$count = 5333;
	#10 counter$count = 5334;
	#10 counter$count = 5335;
	#10 counter$count = 5336;
	#10 counter$count = 5337;
	#10 counter$count = 5338;
	#10 counter$count = 5339;
	#10 counter$count = 5340;
	#10 counter$count = 5341;
	#10 counter$count = 5342;
	#10 counter$count = 5343;
	#10 counter$count = 5344;
	#10 counter$count = 5345;
	#10 counter$count = 5346;
	#10 counter$count = 5347;
	#10 counter$count = 5348;
	#10 counter$count = 5349;
	#10 counter$count = 5350;
	#10 counter$count = 5351;
	#10 counter$count = 5352;
	#10 counter$count = 5353;
	#10 counter$count = 5354;
	#10 counter$count = 5355;
	#10 counter$count = 5356;
	#10 counter$count = 5357;
	#10 counter$count = 5358;
	#10 counter$count = 5359;
	#10 counter$count = 5360;
	#10 counter$count = 5361;
	#10 counter$count = 5362;
	#10 counter$count = 5363;
	#10 counter$count = 5364;
	#10 counter$count = 5365;
	#10 counter$count = 5366;
	#10 counter$count = 5367;
	#10 counter$count = 5368;
	#10 counter$count = 5369;
	#10 counter$count = 5370;
	#10 counter$count = 5371;
	#10 counter$count = 5372;
	#10 counter$count = 5373;
	#10 counter$count = 5374;
	#10 counter$count = 5375;
	#10 counter$count = 5376;
	#10 counter$count = 5377;
	#10 counter$count = 5378;
	#10 counter$count = 5379;
	#10 counter$count = 5380;
	#10 counter$count = 5381;
	#10 counter$count = 5382;
	#10 counter$count = 5383;
	#10 counter$count = 5384;
	#10 counter$count = 5385;
	#10 counter$count = 5386;
	#10 counter$count = 5387;
	#10 counter$count = 5388;
	#10 counter$count = 5389;
	#10 counter$count = 5390;
	#10 counter$count = 5391;
	#10 counter$count = 5392;
	#10 counter$count = 5393;
	#10 counter$count = 5394;
	#10 counter$count = 5395;
	#10 counter$count = 5396;
	#10 counter$count = 5397;
	#10 counter$count = 5398;
	#10 counter$count = 5399;
	#10 counter$count = 5400;
	#10 counter$count = 5401;
	#10 counter$count = 5402;
	#10 counter$count = 5403;
	#10 counter$count = 5404;
	#10 counter$count = 5405;
	#10 counter$count = 5406;
	#10 counter$count = 5407;
	#10 counter$count = 5408;
	#10 counter$count = 5409;
	#10 counter$count = 5410;
	#10 counter$count = 5411;
	#10 counter$count = 5412;
	#10 counter$count = 5413;
	#10 counter$count = 5414;
	#10 counter$count = 5415;
	#10 counter$count = 5416;
	#10 counter$count = 5417;
	#10 counter$count = 5418;
	#10 counter$count = 5419;
	#10 counter$count = 5420;
	#10 counter$count = 5421;
	#10 counter$count = 5422;
	#10 counter$count = 5423;
	#10 counter$count = 5424;
	#10 counter$count = 5425;
	#10 counter$count = 5426;
	#10 counter$count = 5427;
	#10 counter$count = 5428;
	#10 counter$count = 5429;
	#10 counter$count = 5430;
	#10 counter$count = 5431;
	#10 counter$count = 5432;
	#10 counter$count = 5433;
	#10 counter$count = 5434;
	#10 counter$count = 5435;
	#10 counter$count = 5436;
	#10 counter$count = 5437;
	#10 counter$count = 5438;
	#10 counter$count = 5439;
	#10 counter$count = 5440;
	#10 counter$count = 5441;
	#10 counter$count = 5442;
	#10 counter$count = 5443;
	#10 counter$count = 5444;
	#10 counter$count = 5445;
	#10 counter$count = 5446;
	#10 counter$count = 5447;
	#10 counter$count = 5448;
	#10 counter$count = 5449;
	#10 counter$count = 5450;
	#10 counter$count = 5451;
	#10 counter$count = 5452;
	#10 counter$count = 5453;
	#10 counter$count = 5454;
	#10 counter$count = 5455;
	#10 counter$count = 5456;
	#10 counter$count = 5457;
	#10 counter$count = 5458;
	#10 counter$count = 5459;
	#10 counter$count = 5460;
	#10 counter$count = 5461;
	#10 counter$count = 5462;
	#10 counter$count = 5463;
	#10 counter$count = 5464;
	#10 counter$count = 5465;
	#10 counter$count = 5466;
	#10 counter$count = 5467;
	#10 counter$count = 5468;
	#10 counter$count = 5469;
	#10 counter$count = 5470;
	#10 counter$count = 5471;
	#10 counter$count = 5472;
	#10 counter$count = 5473;
	#10 counter$count = 5474;
	#10 counter$count = 5475;
	#10 counter$count = 5476;
	#10 counter$count = 5477;
	#10 counter$count = 5478;
	#10 counter$count = 5479;
	#10 counter$count = 5480;
	#10 counter$count = 5481;
	#10 counter$count = 5482;
	#10 counter$count = 5483;
	#10 counter$count = 5484;
	#10 counter$count = 5485;
	#10 counter$count = 5486;
	#10 counter$count = 5487;
	#10 counter$count = 5488;
	#10 counter$count = 5489;
	#10 counter$count = 5490;
	#10 counter$count = 5491;
	#10 counter$count = 5492;
	#10 counter$count = 5493;
	#10 counter$count = 5494;
	#10 counter$count = 5495;
	#10 counter$count = 5496;
	#10 counter$count = 5497;
	#10 counter$count = 5498;
	#10 counter$count = 5499;
	#10 counter$count = 5500;
	#10 counter$count = 5501;
	#10 counter$count = 5502;
	#10 counter$count = 5503;
	#10 counter$count = 5504;
	#10 counter$count = 5505;
	#10 counter$count = 5506;
	#10 counter$count = 5507;
	#10 counter$count = 5508;
	#10 counter$count = 5509;
	#10 counter$count = 5510;
	#10 counter$count = 5511;
	#10 counter$count = 5512;
	#10 counter$count = 5513;
	#10 counter$count = 5514;
	#10 counter$count = 5515;
	#10 counter$count = 5516;
	#10 counter$count = 5517;
	#10 counter$count = 5518;
	#10 counter$count = 5519;
	#10 counter$count = 5520;
	#10 counter$count = 5521;
	#10 counter$count = 5522;
	#10 counter$count = 5523;
	#10 counter$count = 5524;
	#10 counter$count = 5525;
	#10 counter$count = 5526;
	#10 counter$count = 5527;
	#10 counter$count = 5528;
	#10 counter$count = 5529;
	#10 counter$count = 5530;
	#10 counter$count = 5531;
	#10 counter$count = 5532;
	#10 counter$count = 5533;
	#10 counter$count = 5534;
	#10 counter$count = 5535;
	#10 counter$count = 5536;
	#10 counter$count = 5537;
	#10 counter$count = 5538;
	#10 counter$count = 5539;
	#10 counter$count = 5540;
	#10 counter$count = 5541;
	#10 counter$count = 5542;
	#10 counter$count = 5543;
	#10 counter$count = 5544;
	#10 counter$count = 5545;
	#10 counter$count = 5546;
	#10 counter$count = 5547;
	#10 counter$count = 5548;
	#10 counter$count = 5549;
	#10 counter$count = 5550;
	#10 counter$count = 5551;
	#10 counter$count = 5552;
	#10 counter$count = 5553;
	#10 counter$count = 5554;
	#10 counter$count = 5555;
	#10 counter$count = 5556;
	#10 counter$count = 5557;
	#10 counter$count = 5558;
	#10 counter$count = 5559;
	#10 counter$count = 5560;
	#10 counter$count = 5561;
	#10 counter$count = 5562;
	#10 counter$count = 5563;
	#10 counter$count = 5564;
	#10 counter$count = 5565;
	#10 counter$count = 5566;
	#10 counter$count = 5567;
	#10 counter$count = 5568;
	#10 counter$count = 5569;
	#10 counter$count = 5570;
	#10 counter$count = 5571;
	#10 counter$count = 5572;
	#10 counter$count = 5573;
	#10 counter$count = 5574;
	#10 counter$count = 5575;
	#10 counter$count = 5576;
	#10 counter$count = 5577;
	#10 counter$count = 5578;
	#10 counter$count = 5579;
	#10 counter$count = 5580;
	#10 counter$count = 5581;
	#10 counter$count = 5582;
	#10 counter$count = 5583;
	#10 counter$count = 5584;
	#10 counter$count = 5585;
	#10 counter$count = 5586;
	#10 counter$count = 5587;
	#10 counter$count = 5588;
	#10 counter$count = 5589;
	#10 counter$count = 5590;
	#10 counter$count = 5591;
	#10 counter$count = 5592;
	#10 counter$count = 5593;
	#10 counter$count = 5594;
	#10 counter$count = 5595;
	#10 counter$count = 5596;
	#10 counter$count = 5597;
	#10 counter$count = 5598;
	#10 counter$count = 5599;
	#10 counter$count = 5600;
	#10 counter$count = 5601;
	#10 counter$count = 5602;
	#10 counter$count = 5603;
	#10 counter$count = 5604;
	#10 counter$count = 5605;
	#10 counter$count = 5606;
	#10 counter$count = 5607;
	#10 counter$count = 5608;
	#10 counter$count = 5609;
	#10 counter$count = 5610;
	#10 counter$count = 5611;
	#10 counter$count = 5612;
	#10 counter$count = 5613;
	#10 counter$count = 5614;
	#10 counter$count = 5615;
	#10 counter$count = 5616;
	#10 counter$count = 5617;
	#10 counter$count = 5618;
	#10 counter$count = 5619;
	#10 counter$count = 5620;
	#10 counter$count = 5621;
	#10 counter$count = 5622;
	#10 counter$count = 5623;
	#10 counter$count = 5624;
	#10 counter$count = 5625;
	#10 counter$count = 5626;
	#10 counter$count = 5627;
	#10 counter$count = 5628;
	#10 counter$count = 5629;
	#10 counter$count = 5630;
	#10 counter$count = 5631;
	#10 counter$count = 5632;
	#10 counter$count = 5633;
	#10 counter$count = 5634;
	#10 counter$count = 5635;
	#10 counter$count = 5636;
	#10 counter$count = 5637;
	#10 counter$count = 5638;
	#10 counter$count = 5639;
	#10 counter$count = 5640;
	#10 counter$count = 5641;
	#10 counter$count = 5642;
	#10 counter$count = 5643;
	#10 counter$count = 5644;
	#10 counter$count = 5645;
	#10 counter$count = 5646;
	#10 counter$count = 5647;
	#10 counter$count = 5648;
	#10 counter$count = 5649;
	#10 counter$count = 5650;
	#10 counter$count = 5651;
	#10 counter$count = 5652;
	#10 counter$count = 5653;
	#10 counter$count = 5654;
	#10 counter$count = 5655;
	#10 counter$count = 5656;
	#10 counter$count = 5657;
	#10 counter$count = 5658;
	#10 counter$count = 5659;
	#10 counter$count = 5660;
	#10 counter$count = 5661;
	#10 counter$count = 5662;
	#10 counter$count = 5663;
	#10 counter$count = 5664;
	#10 counter$count = 5665;
	#10 counter$count = 5666;
	#10 counter$count = 5667;
	#10 counter$count = 5668;
	#10 counter$count = 5669;
	#10 counter$count = 5670;
	#10 counter$count = 5671;
	#10 counter$count = 5672;
	#10 counter$count = 5673;
	#10 counter$count = 5674;
	#10 counter$count = 5675;
	#10 counter$count = 5676;
	#10 counter$count = 5677;
	#10 counter$count = 5678;
	#10 counter$count = 5679;
	#10 counter$count = 5680;
	#10 counter$count = 5681;
	#10 counter$count = 5682;
	#10 counter$count = 5683;
	#10 counter$count = 5684;
	#10 counter$count = 5685;
	#10 counter$count = 5686;
	#10 counter$count = 5687;
	#10 counter$count = 5688;
	#10 counter$count = 5689;
	#10 counter$count = 5690;
	#10 counter$count = 5691;
	#10 counter$count = 5692;
	#10 counter$count = 5693;
	#10 counter$count = 5694;
	#10 counter$count = 5695;
	#10 counter$count = 5696;
	#10 counter$count = 5697;
	#10 counter$count = 5698;
	#10 counter$count = 5699;
	#10 counter$count = 5700;
	#10 counter$count = 5701;
	#10 counter$count = 5702;
	#10 counter$count = 5703;
	#10 counter$count = 5704;
	#10 counter$count = 5705;
	#10 counter$count = 5706;
	#10 counter$count = 5707;
	#10 counter$count = 5708;
	#10 counter$count = 5709;
	#10 counter$count = 5710;
	#10 counter$count = 5711;
	#10 counter$count = 5712;
	#10 counter$count = 5713;
	#10 counter$count = 5714;
	#10 counter$count = 5715;
	#10 counter$count = 5716;
	#10 counter$count = 5717;
	#10 counter$count = 5718;
	#10 counter$count = 5719;
	#10 counter$count = 5720;
	#10 counter$count = 5721;
	#10 counter$count = 5722;
	#10 counter$count = 5723;
	#10 counter$count = 5724;
	#10 counter$count = 5725;
	#10 counter$count = 5726;
	#10 counter$count = 5727;
	#10 counter$count = 5728;
	#10 counter$count = 5729;
	#10 counter$count = 5730;
	#10 counter$count = 5731;
	#10 counter$count = 5732;
	#10 counter$count = 5733;
	#10 counter$count = 5734;
	#10 counter$count = 5735;
	#10 counter$count = 5736;
	#10 counter$count = 5737;
	#10 counter$count = 5738;
	#10 counter$count = 5739;
	#10 counter$count = 5740;
	#10 counter$count = 5741;
	#10 counter$count = 5742;
	#10 counter$count = 5743;
	#10 counter$count = 5744;
	#10 counter$count = 5745;
	#10 counter$count = 5746;
	#10 counter$count = 5747;
	#10 counter$count = 5748;
	#10 counter$count = 5749;
	#10 counter$count = 5750;
	#10 counter$count = 5751;
	#10 counter$count = 5752;
	#10 counter$count = 5753;
	#10 counter$count = 5754;
	#10 counter$count = 5755;
	#10 counter$count = 5756;
	#10 counter$count = 5757;
	#10 counter$count = 5758;
	#10 counter$count = 5759;
	#10 counter$count = 5760;
	#10 counter$count = 5761;
	#10 counter$count = 5762;
	#10 counter$count = 5763;
	#10 counter$count = 5764;
	#10 counter$count = 5765;
	#10 counter$count = 5766;
	#10 counter$count = 5767;
	#10 counter$count = 5768;
	#10 counter$count = 5769;
	#10 counter$count = 5770;
	#10 counter$count = 5771;
	#10 counter$count = 5772;
	#10 counter$count = 5773;
	#10 counter$count = 5774;
	#10 counter$count = 5775;
	#10 counter$count = 5776;
	#10 counter$count = 5777;
	#10 counter$count = 5778;
	#10 counter$count = 5779;
	#10 counter$count = 5780;
	#10 counter$count = 5781;
	#10 counter$count = 5782;
	#10 counter$count = 5783;
	#10 counter$count = 5784;
	#10 counter$count = 5785;
	#10 counter$count = 5786;
	#10 counter$count = 5787;
	#10 counter$count = 5788;
	#10 counter$count = 5789;
	#10 counter$count = 5790;
	#10 counter$count = 5791;
	#10 counter$count = 5792;
	#10 counter$count = 5793;
	#10 counter$count = 5794;
	#10 counter$count = 5795;
	#10 counter$count = 5796;
	#10 counter$count = 5797;
	#10 counter$count = 5798;
	#10 counter$count = 5799;
	#10 counter$count = 5800;
	#10 counter$count = 5801;
	#10 counter$count = 5802;
	#10 counter$count = 5803;
	#10 counter$count = 5804;
	#10 counter$count = 5805;
	#10 counter$count = 5806;
	#10 counter$count = 5807;
	#10 counter$count = 5808;
	#10 counter$count = 5809;
	#10 counter$count = 5810;
	#10 counter$count = 5811;
	#10 counter$count = 5812;
	#10 counter$count = 5813;
	#10 counter$count = 5814;
	#10 counter$count = 5815;
	#10 counter$count = 5816;
	#10 counter$count = 5817;
	#10 counter$count = 5818;
	#10 counter$count = 5819;
	#10 counter$count = 5820;
	#10 counter$count = 5821;
	#10 counter$count = 5822;
	#10 counter$count = 5823;
	#10 counter$count = 5824;
	#10 counter$count = 5825;
	#10 counter$count = 5826;
	#10 counter$count = 5827;
	#10 counter$count = 5828;
	#10 counter$count = 5829;
	#10 counter$count = 5830;
	#10 counter$count = 5831;
	#10 counter$count = 5832;
	#10 counter$count = 5833;
	#10 counter$count = 5834;
	#10 counter$count = 5835;
	#10 counter$count = 5836;
	#10 counter$count = 5837;
	#10 counter$count = 5838;
	#10 counter$count = 5839;
	#10 counter$count = 5840;
	#10 counter$count = 5841;
	#10 counter$count = 5842;
	#10 counter$count = 5843;
	#10 counter$count = 5844;
	#10 counter$count = 5845;
	#10 counter$count = 5846;
	#10 counter$count = 5847;
	#10 counter$count = 5848;
	#10 counter$count = 5849;
	#10 counter$count = 5850;
	#10 counter$count = 5851;
	#10 counter$count = 5852;
	#10 counter$count = 5853;
	#10 counter$count = 5854;
	#10 counter$count = 5855;
	#10 counter$count = 5856;
	#10 counter$count = 5857;
	#10 counter$count = 5858;
	#10 counter$count = 5859;
	#10 counter$count = 5860;
	#10 counter$count = 5861;
	#10 counter$count = 5862;
	#10 counter$count = 5863;
	#10 counter$count = 5864;
	#10 counter$count = 5865;
	#10 counter$count = 5866;
	#10 counter$count = 5867;
	#10 counter$count = 5868;
	#10 counter$count = 5869;
	#10 counter$count = 5870;
	#10 counter$count = 5871;
	#10 counter$count = 5872;
	#10 counter$count = 5873;
	#10 counter$count = 5874;
	#10 counter$count = 5875;
	#10 counter$count = 5876;
	#10 counter$count = 5877;
	#10 counter$count = 5878;
	#10 counter$count = 5879;
	#10 counter$count = 5880;
	#10 counter$count = 5881;
	#10 counter$count = 5882;
	#10 counter$count = 5883;
	#10 counter$count = 5884;
	#10 counter$count = 5885;
	#10 counter$count = 5886;
	#10 counter$count = 5887;
	#10 counter$count = 5888;
	#10 counter$count = 5889;
	#10 counter$count = 5890;
	#10 counter$count = 5891;
	#10 counter$count = 5892;
	#10 counter$count = 5893;
	#10 counter$count = 5894;
	#10 counter$count = 5895;
	#10 counter$count = 5896;
	#10 counter$count = 5897;
	#10 counter$count = 5898;
	#10 counter$count = 5899;
	#10 counter$count = 5900;
	#10 counter$count = 5901;
	#10 counter$count = 5902;
	#10 counter$count = 5903;
	#10 counter$count = 5904;
	#10 counter$count = 5905;
	#10 counter$count = 5906;
	#10 counter$count = 5907;
	#10 counter$count = 5908;
	#10 counter$count = 5909;
	#10 counter$count = 5910;
	#10 counter$count = 5911;
	#10 counter$count = 5912;
	#10 counter$count = 5913;
	#10 counter$count = 5914;
	#10 counter$count = 5915;
	#10 counter$count = 5916;
	#10 counter$count = 5917;
	#10 counter$count = 5918;
	#10 counter$count = 5919;
	#10 counter$count = 5920;
	#10 counter$count = 5921;
	#10 counter$count = 5922;
	#10 counter$count = 5923;
	#10 counter$count = 5924;
	#10 counter$count = 5925;
	#10 counter$count = 5926;
	#10 counter$count = 5927;
	#10 counter$count = 5928;
	#10 counter$count = 5929;
	#10 counter$count = 5930;
	#10 counter$count = 5931;
	#10 counter$count = 5932;
	#10 counter$count = 5933;
	#10 counter$count = 5934;
	#10 counter$count = 5935;
	#10 counter$count = 5936;
	#10 counter$count = 5937;
	#10 counter$count = 5938;
	#10 counter$count = 5939;
	#10 counter$count = 5940;
	#10 counter$count = 5941;
	#10 counter$count = 5942;
	#10 counter$count = 5943;
	#10 counter$count = 5944;
	#10 counter$count = 5945;
	#10 counter$count = 5946;
	#10 counter$count = 5947;
	#10 counter$count = 5948;
	#10 counter$count = 5949;
	#10 counter$count = 5950;
	#10 counter$count = 5951;
	#10 counter$count = 5952;
	#10 counter$count = 5953;
	#10 counter$count = 5954;
	#10 counter$count = 5955;
	#10 counter$count = 5956;
	#10 counter$count = 5957;
	#10 counter$count = 5958;
	#10 counter$count = 5959;
	#10 counter$count = 5960;
	#10 counter$count = 5961;
	#10 counter$count = 5962;
	#10 counter$count = 5963;
	#10 counter$count = 5964;
	#10 counter$count = 5965;
	#10 counter$count = 5966;
	#10 counter$count = 5967;
	#10 counter$count = 5968;
	#10 counter$count = 5969;
	#10 counter$count = 5970;
	#10 counter$count = 5971;
	#10 counter$count = 5972;
	#10 counter$count = 5973;
	#10 counter$count = 5974;
	#10 counter$count = 5975;
	#10 counter$count = 5976;
	#10 counter$count = 5977;
	#10 counter$count = 5978;
	#10 counter$count = 5979;
	#10 counter$count = 5980;
	#10 counter$count = 5981;
	#10 counter$count = 5982;
	#10 counter$count = 5983;
	#10 counter$count = 5984;
	#10 counter$count = 5985;
	#10 counter$count = 5986;
	#10 counter$count = 5987;
	#10 counter$count = 5988;
	#10 counter$count = 5989;
	#10 counter$count = 5990;
	#10 counter$count = 5991;
	#10 counter$count = 5992;
	#10 counter$count = 5993;
	#10 counter$count = 5994;
	#10 counter$count = 5995;
	#10 counter$count = 5996;
	#10 counter$count = 5997;
	#10 counter$count = 5998;
	#10 counter$count = 5999;
	#10 counter$count = 6000;
	#10 counter$count = 6001;
	#10 counter$count = 6002;
	#10 counter$count = 6003;
	#10 counter$count = 6004;
	#10 counter$count = 6005;
	#10 counter$count = 6006;
	#10 counter$count = 6007;
	#10 counter$count = 6008;
	#10 counter$count = 6009;
	#10 counter$count = 6010;
	#10 counter$count = 6011;
	#10 counter$count = 6012;
	#10 counter$count = 6013;
	#10 counter$count = 6014;
	#10 counter$count = 6015;
	#10 counter$count = 6016;
	#10 counter$count = 6017;
	#10 counter$count = 6018;
	#10 counter$count = 6019;
	#10 counter$count = 6020;
	#10 counter$count = 6021;
	#10 counter$count = 6022;
	#10 counter$count = 6023;
	#10 counter$count = 6024;
	#10 counter$count = 6025;
	#10 counter$count = 6026;
	#10 counter$count = 6027;
	#10 counter$count = 6028;
	#10 counter$count = 6029;
	#10 counter$count = 6030;
	#10 counter$count = 6031;
	#10 counter$count = 6032;
	#10 counter$count = 6033;
	#10 counter$count = 6034;
	#10 counter$count = 6035;
	#10 counter$count = 6036;
	#10 counter$count = 6037;
	#10 counter$count = 6038;
	#10 counter$count = 6039;
	#10 counter$count = 6040;
	#10 counter$count = 6041;
	#10 counter$count = 6042;
	#10 counter$count = 6043;
	#10 counter$count = 6044;
	#10 counter$count = 6045;
	#10 counter$count = 6046;
	#10 counter$count = 6047;
	#10 counter$count = 6048;
	#10 counter$count = 6049;
	#10 counter$count = 6050;
	#10 counter$count = 6051;
	#10 counter$count = 6052;
	#10 counter$count = 6053;
	#10 counter$count = 6054;
	#10 counter$count = 6055;
	#10 counter$count = 6056;
	#10 counter$count = 6057;
	#10 counter$count = 6058;
	#10 counter$count = 6059;
	#10 counter$count = 6060;
	#10 counter$count = 6061;
	#10 counter$count = 6062;
	#10 counter$count = 6063;
	#10 counter$count = 6064;
	#10 counter$count = 6065;
	#10 counter$count = 6066;
	#10 counter$count = 6067;
	#10 counter$count = 6068;
	#10 counter$count = 6069;
	#10 counter$count = 6070;
	#10 counter$count = 6071;
	#10 counter$count = 6072;
	#10 counter$count = 6073;
	#10 counter$count = 6074;
	#10 counter$count = 6075;
	#10 counter$count = 6076;
	#10 counter$count = 6077;
	#10 counter$count = 6078;
	#10 counter$count = 6079;
	#10 counter$count = 6080;
	#10 counter$count = 6081;
	#10 counter$count = 6082;
	#10 counter$count = 6083;
	#10 counter$count = 6084;
	#10 counter$count = 6085;
	#10 counter$count = 6086;
	#10 counter$count = 6087;
	#10 counter$count = 6088;
	#10 counter$count = 6089;
	#10 counter$count = 6090;
	#10 counter$count = 6091;
	#10 counter$count = 6092;
	#10 counter$count = 6093;
	#10 counter$count = 6094;
	#10 counter$count = 6095;
	#10 counter$count = 6096;
	#10 counter$count = 6097;
	#10 counter$count = 6098;
	#10 counter$count = 6099;
	#10 counter$count = 6100;
	#10 counter$count = 6101;
	#10 counter$count = 6102;
	#10 counter$count = 6103;
	#10 counter$count = 6104;
	#10 counter$count = 6105;
	#10 counter$count = 6106;
	#10 counter$count = 6107;
	#10 counter$count = 6108;
	#10 counter$count = 6109;
	#10 counter$count = 6110;
	#10 counter$count = 6111;
	#10 counter$count = 6112;
	#10 counter$count = 6113;
	#10 counter$count = 6114;
	#10 counter$count = 6115;
	#10 counter$count = 6116;
	#10 counter$count = 6117;
	#10 counter$count = 6118;
	#10 counter$count = 6119;
	#10 counter$count = 6120;
	#10 counter$count = 6121;
	#10 counter$count = 6122;
	#10 counter$count = 6123;
	#10 counter$count = 6124;
	#10 counter$count = 6125;
	#10 counter$count = 6126;
	#10 counter$count = 6127;
	#10 counter$count = 6128;
	#10 counter$count = 6129;
	#10 counter$count = 6130;
	#10 counter$count = 6131;
	#10 counter$count = 6132;
	#10 counter$count = 6133;
	#10 counter$count = 6134;
	#10 counter$count = 6135;
	#10 counter$count = 6136;
	#10 counter$count = 6137;
	#10 counter$count = 6138;
	#10 counter$count = 6139;
	#10 counter$count = 6140;
	#10 counter$count = 6141;
	#10 counter$count = 6142;
	#10 counter$count = 6143;
	#10 counter$count = 6144;
	#10 counter$count = 6145;
	#10 counter$count = 6146;
	#10 counter$count = 6147;
	#10 counter$count = 6148;
	#10 counter$count = 6149;
	#10 counter$count = 6150;
	#10 counter$count = 6151;
	#10 counter$count = 6152;
	#10 counter$count = 6153;
	#10 counter$count = 6154;
	#10 counter$count = 6155;
	#10 counter$count = 6156;
	#10 counter$count = 6157;
	#10 counter$count = 6158;
	#10 counter$count = 6159;
	#10 counter$count = 6160;
	#10 counter$count = 6161;
	#10 counter$count = 6162;
	#10 counter$count = 6163;
	#10 counter$count = 6164;
	#10 counter$count = 6165;
	#10 counter$count = 6166;
	#10 counter$count = 6167;
	#10 counter$count = 6168;
	#10 counter$count = 6169;
	#10 counter$count = 6170;
	#10 counter$count = 6171;
	#10 counter$count = 6172;
	#10 counter$count = 6173;
	#10 counter$count = 6174;
	#10 counter$count = 6175;
	#10 counter$count = 6176;
	#10 counter$count = 6177;
	#10 counter$count = 6178;
	#10 counter$count = 6179;
	#10 counter$count = 6180;
	#10 counter$count = 6181;
	#10 counter$count = 6182;
	#10 counter$count = 6183;
	#10 counter$count = 6184;
	#10 counter$count = 6185;
	#10 counter$count = 6186;
	#10 counter$count = 6187;
	#10 counter$count = 6188;
	#10 counter$count = 6189;
	#10 counter$count = 6190;
	#10 counter$count = 6191;
	#10 counter$count = 6192;
	#10 counter$count = 6193;
	#10 counter$count = 6194;
	#10 counter$count = 6195;
	#10 counter$count = 6196;
	#10 counter$count = 6197;
	#10 counter$count = 6198;
	#10 counter$count = 6199;
	#10 counter$count = 6200;
	#10 counter$count = 6201;
	#10 counter$count = 6202;
	#10 counter$count = 6203;
	#10 counter$count = 6204;
	#10 counter$count = 6205;
	#10 counter$count = 6206;
	#10 counter$count = 6207;
	#10 counter$count = 6208;
	#10 counter$count = 6209;
	#10 counter$count = 6210;
	#10 counter$count = 6211;
	#10 counter$count = 6212;
	#10 counter$count = 6213;
	#10 counter$count = 6214;
	#10 counter$count = 6215;
	#10 counter$count = 6216;
	#10 counter$count = 6217;
	#10 counter$count = 6218;
	#10 counter$count = 6219;
	#10 counter$count = 6220;
	#10 counter$count = 6221;
	#10 counter$count = 6222;
	#10 counter$count = 6223;
	#10 counter$count = 6224;
	#10 counter$count = 6225;
	#10 counter$count = 6226;
	#10 counter$count = 6227;
	#10 counter$count = 6228;
	#10 counter$count = 6229;
	#10 counter$count = 6230;
	#10 counter$count = 6231;
	#10 counter$count = 6232;
	#10 counter$count = 6233;
	#10 counter$count = 6234;
	#10 counter$count = 6235;
	#10 counter$count = 6236;
	#10 counter$count = 6237;
	#10 counter$count = 6238;
	#10 counter$count = 6239;
	#10 counter$count = 6240;
	#10 counter$count = 6241;
	#10 counter$count = 6242;
	#10 counter$count = 6243;
	#10 counter$count = 6244;
	#10 counter$count = 6245;
	#10 counter$count = 6246;
	#10 counter$count = 6247;
	#10 counter$count = 6248;
	#10 counter$count = 6249;
	#10 counter$count = 6250;
	#10 counter$count = 6251;
	#10 counter$count = 6252;
	#10 counter$count = 6253;
	#10 counter$count = 6254;
	#10 counter$count = 6255;
	#10 counter$count = 6256;
	#10 counter$count = 6257;
	#10 counter$count = 6258;
	#10 counter$count = 6259;
	#10 counter$count = 6260;
	#10 counter$count = 6261;
	#10 counter$count = 6262;
	#10 counter$count = 6263;
	#10 counter$count = 6264;
	#10 counter$count = 6265;
	#10 counter$count = 6266;
	#10 counter$count = 6267;
	#10 counter$count = 6268;
	#10 counter$count = 6269;
	#10 counter$count = 6270;
	#10 counter$count = 6271;
	#10 counter$count = 6272;
	#10 counter$count = 6273;
	#10 counter$count = 6274;
	#10 counter$count = 6275;
	#10 counter$count = 6276;
	#10 counter$count = 6277;
	#10 counter$count = 6278;
	#10 counter$count = 6279;
	#10 counter$count = 6280;
	#10 counter$count = 6281;
	#10 counter$count = 6282;
	#10 counter$count = 6283;
	#10 counter$count = 6284;
	#10 counter$count = 6285;
	#10 counter$count = 6286;
	#10 counter$count = 6287;
	#10 counter$count = 6288;
	#10 counter$count = 6289;
	#10 counter$count = 6290;
	#10 counter$count = 6291;
	#10 counter$count = 6292;
	#10 counter$count = 6293;
	#10 counter$count = 6294;
	#10 counter$count = 6295;
	#10 counter$count = 6296;
	#10 counter$count = 6297;
	#10 counter$count = 6298;
	#10 counter$count = 6299;
	#10 counter$count = 6300;
	#10 counter$count = 6301;
	#10 counter$count = 6302;
	#10 counter$count = 6303;
	#10 counter$count = 6304;
	#10 counter$count = 6305;
	#10 counter$count = 6306;
	#10 counter$count = 6307;
	#10 counter$count = 6308;
	#10 counter$count = 6309;
	#10 counter$count = 6310;
	#10 counter$count = 6311;
	#10 counter$count = 6312;
	#10 counter$count = 6313;
	#10 counter$count = 6314;
	#10 counter$count = 6315;
	#10 counter$count = 6316;
	#10 counter$count = 6317;
	#10 counter$count = 6318;
	#10 counter$count = 6319;
	#10 counter$count = 6320;
	#10 counter$count = 6321;
	#10 counter$count = 6322;
	#10 counter$count = 6323;
	#10 counter$count = 6324;
	#10 counter$count = 6325;
	#10 counter$count = 6326;
	#10 counter$count = 6327;
	#10 counter$count = 6328;
	#10 counter$count = 6329;
	#10 counter$count = 6330;
	#10 counter$count = 6331;
	#10 counter$count = 6332;
	#10 counter$count = 6333;
	#10 counter$count = 6334;
	#10 counter$count = 6335;
	#10 counter$count = 6336;
	#10 counter$count = 6337;
	#10 counter$count = 6338;
	#10 counter$count = 6339;
	#10 counter$count = 6340;
	#10 counter$count = 6341;
	#10 counter$count = 6342;
	#10 counter$count = 6343;
	#10 counter$count = 6344;
	#10 counter$count = 6345;
	#10 counter$count = 6346;
	#10 counter$count = 6347;
	#10 counter$count = 6348;
	#10 counter$count = 6349;
	#10 counter$count = 6350;
	#10 counter$count = 6351;
	#10 counter$count = 6352;
	#10 counter$count = 6353;
	#10 counter$count = 6354;
	#10 counter$count = 6355;
	#10 counter$count = 6356;
	#10 counter$count = 6357;
	#10 counter$count = 6358;
	#10 counter$count = 6359;
	#10 counter$count = 6360;
	#10 counter$count = 6361;
	#10 counter$count = 6362;
	#10 counter$count = 6363;
	#10 counter$count = 6364;
	#10 counter$count = 6365;
	#10 counter$count = 6366;
	#10 counter$count = 6367;
	#10 counter$count = 6368;
	#10 counter$count = 6369;
	#10 counter$count = 6370;
	#10 counter$count = 6371;
	#10 counter$count = 6372;
	#10 counter$count = 6373;
	#10 counter$count = 6374;
	#10 counter$count = 6375;
	#10 counter$count = 6376;
	#10 counter$count = 6377;
	#10 counter$count = 6378;
	#10 counter$count = 6379;
	#10 counter$count = 6380;
	#10 counter$count = 6381;
	#10 counter$count = 6382;
	#10 counter$count = 6383;
	#10 counter$count = 6384;
	#10 counter$count = 6385;
	#10 counter$count = 6386;
	#10 counter$count = 6387;
	#10 counter$count = 6388;
	#10 counter$count = 6389;
	#10 counter$count = 6390;
	#10 counter$count = 6391;
	#10 counter$count = 6392;
	#10 counter$count = 6393;
	#10 counter$count = 6394;
	#10 counter$count = 6395;
	#10 counter$count = 6396;
	#10 counter$count = 6397;
	#10 counter$count = 6398;
	#10 counter$count = 6399;
	#10 counter$count = 6400;
	#10 counter$count = 6401;
	#10 counter$count = 6402;
	#10 counter$count = 6403;
	#10 counter$count = 6404;
	#10 counter$count = 6405;
	#10 counter$count = 6406;
	#10 counter$count = 6407;
	#10 counter$count = 6408;
	#10 counter$count = 6409;
	#10 counter$count = 6410;
	#10 counter$count = 6411;
	#10 counter$count = 6412;
	#10 counter$count = 6413;
	#10 counter$count = 6414;
	#10 counter$count = 6415;
	#10 counter$count = 6416;
	#10 counter$count = 6417;
	#10 counter$count = 6418;
	#10 counter$count = 6419;
	#10 counter$count = 6420;
	#10 counter$count = 6421;
	#10 counter$count = 6422;
	#10 counter$count = 6423;
	#10 counter$count = 6424;
	#10 counter$count = 6425;
	#10 counter$count = 6426;
	#10 counter$count = 6427;
	#10 counter$count = 6428;
	#10 counter$count = 6429;
	#10 counter$count = 6430;
	#10 counter$count = 6431;
	#10 counter$count = 6432;
	#10 counter$count = 6433;
	#10 counter$count = 6434;
	#10 counter$count = 6435;
	#10 counter$count = 6436;
	#10 counter$count = 6437;
	#10 counter$count = 6438;
	#10 counter$count = 6439;
	#10 counter$count = 6440;
	#10 counter$count = 6441;
	#10 counter$count = 6442;
	#10 counter$count = 6443;
	#10 counter$count = 6444;
	#10 counter$count = 6445;
	#10 counter$count = 6446;
	#10 counter$count = 6447;
	#10 counter$count = 6448;
	#10 counter$count = 6449;
	#10 counter$count = 6450;
	#10 counter$count = 6451;
	#10 counter$count = 6452;
	#10 counter$count = 6453;
	#10 counter$count = 6454;
	#10 counter$count = 6455;
	#10 counter$count = 6456;
	#10 counter$count = 6457;
	#10 counter$count = 6458;
	#10 counter$count = 6459;
	#10 counter$count = 6460;
	#10 counter$count = 6461;
	#10 counter$count = 6462;
	#10 counter$count = 6463;
	#10 counter$count = 6464;
	#10 counter$count = 6465;
	#10 counter$count = 6466;
	#10 counter$count = 6467;
	#10 counter$count = 6468;
	#10 counter$count = 6469;
	#10 counter$count = 6470;
	#10 counter$count = 6471;
	#10 counter$count = 6472;
	#10 counter$count = 6473;
	#10 counter$count = 6474;
	#10 counter$count = 6475;
	#10 counter$count = 6476;
	#10 counter$count = 6477;
	#10 counter$count = 6478;
	#10 counter$count = 6479;
	#10 counter$count = 6480;
	#10 counter$count = 6481;
	#10 counter$count = 6482;
	#10 counter$count = 6483;
	#10 counter$count = 6484;
	#10 counter$count = 6485;
	#10 counter$count = 6486;
	#10 counter$count = 6487;
	#10 counter$count = 6488;
	#10 counter$count = 6489;
	#10 counter$count = 6490;
	#10 counter$count = 6491;
	#10 counter$count = 6492;
	#10 counter$count = 6493;
	#10 counter$count = 6494;
	#10 counter$count = 6495;
	#10 counter$count = 6496;
	#10 counter$count = 6497;
	#10 counter$count = 6498;
	#10 counter$count = 6499;
	#10 counter$count = 6500;
	#10 counter$count = 6501;
	#10 counter$count = 6502;
	#10 counter$count = 6503;
	#10 counter$count = 6504;
	#10 counter$count = 6505;
	#10 counter$count = 6506;
	#10 counter$count = 6507;
	#10 counter$count = 6508;
	#10 counter$count = 6509;
	#10 counter$count = 6510;
	#10 counter$count = 6511;
	#10 counter$count = 6512;
	#10 counter$count = 6513;
	#10 counter$count = 6514;
	#10 counter$count = 6515;
	#10 counter$count = 6516;
	#10 counter$count = 6517;
	#10 counter$count = 6518;
	#10 counter$count = 6519;
	#10 counter$count = 6520;
	#10 counter$count = 6521;
	#10 counter$count = 6522;
	#10 counter$count = 6523;
	#10 counter$count = 6524;
	#10 counter$count = 6525;
	#10 counter$count = 6526;
	#10 counter$count = 6527;
	#10 counter$count = 6528;
	#10 counter$count = 6529;
	#10 counter$count = 6530;
	#10 counter$count = 6531;
	#10 counter$count = 6532;
	#10 counter$count = 6533;
	#10 counter$count = 6534;
	#10 counter$count = 6535;
	#10 counter$count = 6536;
	#10 counter$count = 6537;
	#10 counter$count = 6538;
	#10 counter$count = 6539;
	#10 counter$count = 6540;
	#10 counter$count = 6541;
	#10 counter$count = 6542;
	#10 counter$count = 6543;
	#10 counter$count = 6544;
	#10 counter$count = 6545;
	#10 counter$count = 6546;
	#10 counter$count = 6547;
	#10 counter$count = 6548;
	#10 counter$count = 6549;
	#10 counter$count = 6550;
	#10 counter$count = 6551;
	#10 counter$count = 6552;
	#10 counter$count = 6553;
	#10 counter$count = 6554;
	#10 counter$count = 6555;
	#10 counter$count = 6556;
	#10 counter$count = 6557;
	#10 counter$count = 6558;
	#10 counter$count = 6559;
	#10 counter$count = 6560;
	#10 counter$count = 6561;
	#10 counter$count = 6562;
	#10 counter$count = 6563;
	#10 counter$count = 6564;
	#10 counter$count = 6565;
	#10 counter$count = 6566;
	#10 counter$count = 6567;
	#10 counter$count = 6568;
	#10 counter$count = 6569;
	#10 counter$count = 6570;
	#10 counter$count = 6571;
	#10 counter$count = 6572;
	#10 counter$count = 6573;
	#10 counter$count = 6574;
	#10 counter$count = 6575;
	#10 counter$count = 6576;
	#10 counter$count = 6577;
	#10 counter$count = 6578;
	#10 counter$count = 6579;
	#10 counter$count = 6580;
	#10 counter$count = 6581;
	#10 counter$count = 6582;
	#10 counter$count = 6583;
	#10 counter$count = 6584;
	#10 counter$count = 6585;
	#10 counter$count = 6586;
	#10 counter$count = 6587;
	#10 counter$count = 6588;
	#10 counter$count = 6589;
	#10 counter$count = 6590;
	#10 counter$count = 6591;
	#10 counter$count = 6592;
	#10 counter$count = 6593;
	#10 counter$count = 6594;
	#10 counter$count = 6595;
	#10 counter$count = 6596;
	#10 counter$count = 6597;
	#10 counter$count = 6598;
	#10 counter$count = 6599;
	#10 counter$count = 6600;
	#10 counter$count = 6601;
	#10 counter$count = 6602;
	#10 counter$count = 6603;
	#10 counter$count = 6604;
	#10 counter$count = 6605;
	#10 counter$count = 6606;
	#10 counter$count = 6607;
	#10 counter$count = 6608;
	#10 counter$count = 6609;
	#10 counter$count = 6610;
	#10 counter$count = 6611;
	#10 counter$count = 6612;
	#10 counter$count = 6613;
	#10 counter$count = 6614;
	#10 counter$count = 6615;
	#10 counter$count = 6616;
	#10 counter$count = 6617;
	#10 counter$count = 6618;
	#10 counter$count = 6619;
	#10 counter$count = 6620;
	#10 counter$count = 6621;
	#10 counter$count = 6622;
	#10 counter$count = 6623;
	#10 counter$count = 6624;
	#10 counter$count = 6625;
	#10 counter$count = 6626;
	#10 counter$count = 6627;
	#10 counter$count = 6628;
	#10 counter$count = 6629;
	#10 counter$count = 6630;
	#10 counter$count = 6631;
	#10 counter$count = 6632;
	#10 counter$count = 6633;
	#10 counter$count = 6634;
	#10 counter$count = 6635;
	#10 counter$count = 6636;
	#10 counter$count = 6637;
	#10 counter$count = 6638;
	#10 counter$count = 6639;
	#10 counter$count = 6640;
	#10 counter$count = 6641;
	#10 counter$count = 6642;
	#10 counter$count = 6643;
	#10 counter$count = 6644;
	#10 counter$count = 6645;
	#10 counter$count = 6646;
	#10 counter$count = 6647;
	#10 counter$count = 6648;
	#10 counter$count = 6649;
	#10 counter$count = 6650;
	#10 counter$count = 6651;
	#10 counter$count = 6652;
	#10 counter$count = 6653;
	#10 counter$count = 6654;
	#10 counter$count = 6655;
	#10 counter$count = 6656;
	#10 counter$count = 6657;
	#10 counter$count = 6658;
	#10 counter$count = 6659;
	#10 counter$count = 6660;
	#10 counter$count = 6661;
	#10 counter$count = 6662;
	#10 counter$count = 6663;
	#10 counter$count = 6664;
	#10 counter$count = 6665;
	#10 counter$count = 6666;
	#10 counter$count = 6667;
	#10 counter$count = 6668;
	#10 counter$count = 6669;
	#10 counter$count = 6670;
	#10 counter$count = 6671;
	#10 counter$count = 6672;
	#10 counter$count = 6673;
	#10 counter$count = 6674;
	#10 counter$count = 6675;
	#10 counter$count = 6676;
	#10 counter$count = 6677;
	#10 counter$count = 6678;
	#10 counter$count = 6679;
	#10 counter$count = 6680;
	#10 counter$count = 6681;
	#10 counter$count = 6682;
	#10 counter$count = 6683;
	#10 counter$count = 6684;
	#10 counter$count = 6685;
	#10 counter$count = 6686;
	#10 counter$count = 6687;
	#10 counter$count = 6688;
	#10 counter$count = 6689;
	#10 counter$count = 6690;
	#10 counter$count = 6691;
	#10 counter$count = 6692;
	#10 counter$count = 6693;
	#10 counter$count = 6694;
	#10 counter$count = 6695;
	#10 counter$count = 6696;
	#10 counter$count = 6697;
	#10 counter$count = 6698;
	#10 counter$count = 6699;
	#10 counter$count = 6700;
	#10 counter$count = 6701;
	#10 counter$count = 6702;
	#10 counter$count = 6703;
	#10 counter$count = 6704;
	#10 counter$count = 6705;
	#10 counter$count = 6706;
	#10 counter$count = 6707;
	#10 counter$count = 6708;
	#10 counter$count = 6709;
	#10 counter$count = 6710;
	#10 counter$count = 6711;
	#10 counter$count = 6712;
	#10 counter$count = 6713;
	#10 counter$count = 6714;
	#10 counter$count = 6715;
	#10 counter$count = 6716;
	#10 counter$count = 6717;
	#10 counter$count = 6718;
	#10 counter$count = 6719;
	#10 counter$count = 6720;
	#10 counter$count = 6721;
	#10 counter$count = 6722;
	#10 counter$count = 6723;
	#10 counter$count = 6724;
	#10 counter$count = 6725;
	#10 counter$count = 6726;
	#10 counter$count = 6727;
	#10 counter$count = 6728;
	#10 counter$count = 6729;
	#10 counter$count = 6730;
	#10 counter$count = 6731;
	#10 counter$count = 6732;
	#10 counter$count = 6733;
	#10 counter$count = 6734;
	#10 counter$count = 6735;
	#10 counter$count = 6736;
	#10 counter$count = 6737;
	#10 counter$count = 6738;
	#10 counter$count = 6739;
	#10 counter$count = 6740;
	#10 counter$count = 6741;
	#10 counter$count = 6742;
	#10 counter$count = 6743;
	#10 counter$count = 6744;
	#10 counter$count = 6745;
	#10 counter$count = 6746;
	#10 counter$count = 6747;
	#10 counter$count = 6748;
	#10 counter$count = 6749;
	#10 counter$count = 6750;
	#10 counter$count = 6751;
	#10 counter$count = 6752;
	#10 counter$count = 6753;
	#10 counter$count = 6754;
	#10 counter$count = 6755;
	#10 counter$count = 6756;
	#10 counter$count = 6757;
	#10 counter$count = 6758;
	#10 counter$count = 6759;
	#10 counter$count = 6760;
	#10 counter$count = 6761;
	#10 counter$count = 6762;
	#10 counter$count = 6763;
	#10 counter$count = 6764;
	#10 counter$count = 6765;
	#10 counter$count = 6766;
	#10 counter$count = 6767;
	#10 counter$count = 6768;
	#10 counter$count = 6769;
	#10 counter$count = 6770;
	#10 counter$count = 6771;
	#10 counter$count = 6772;
	#10 counter$count = 6773;
	#10 counter$count = 6774;
	#10 counter$count = 6775;
	#10 counter$count = 6776;
	#10 counter$count = 6777;
	#10 counter$count = 6778;
	#10 counter$count = 6779;
	#10 counter$count = 6780;
	#10 counter$count = 6781;
	#10 counter$count = 6782;
	#10 counter$count = 6783;
	#10 counter$count = 6784;
	#10 counter$count = 6785;
	#10 counter$count = 6786;
	#10 counter$count = 6787;
	#10 counter$count = 6788;
	#10 counter$count = 6789;
	#10 counter$count = 6790;
	#10 counter$count = 6791;
	#10 counter$count = 6792;
	#10 counter$count = 6793;
	#10 counter$count = 6794;
	#10 counter$count = 6795;
	#10 counter$count = 6796;
	#10 counter$count = 6797;
	#10 counter$count = 6798;
	#10 counter$count = 6799;
	#10 counter$count = 6800;
	#10 counter$count = 6801;
	#10 counter$count = 6802;
	#10 counter$count = 6803;
	#10 counter$count = 6804;
	#10 counter$count = 6805;
	#10 counter$count = 6806;
	#10 counter$count = 6807;
	#10 counter$count = 6808;
	#10 counter$count = 6809;
	#10 counter$count = 6810;
	#10 counter$count = 6811;
	#10 counter$count = 6812;
	#10 counter$count = 6813;
	#10 counter$count = 6814;
	#10 counter$count = 6815;
	#10 counter$count = 6816;
	#10 counter$count = 6817;
	#10 counter$count = 6818;
	#10 counter$count = 6819;
	#10 counter$count = 6820;
	#10 counter$count = 6821;
	#10 counter$count = 6822;
	#10 counter$count = 6823;
	#10 counter$count = 6824;
	#10 counter$count = 6825;
	#10 counter$count = 6826;
	#10 counter$count = 6827;
	#10 counter$count = 6828;
	#10 counter$count = 6829;
	#10 counter$count = 6830;
	#10 counter$count = 6831;
	#10 counter$count = 6832;
	#10 counter$count = 6833;
	#10 counter$count = 6834;
	#10 counter$count = 6835;
	#10 counter$count = 6836;
	#10 counter$count = 6837;
	#10 counter$count = 6838;
	#10 counter$count = 6839;
	#10 counter$count = 6840;
	#10 counter$count = 6841;
	#10 counter$count = 6842;
	#10 counter$count = 6843;
	#10 counter$count = 6844;
	#10 counter$count = 6845;
	#10 counter$count = 6846;
	#10 counter$count = 6847;
	#10 counter$count = 6848;
	#10 counter$count = 6849;
	#10 counter$count = 6850;
	#10 counter$count = 6851;
	#10 counter$count = 6852;
	#10 counter$count = 6853;
	#10 counter$count = 6854;
	#10 counter$count = 6855;
	#10 counter$count = 6856;
	#10 counter$count = 6857;
	#10 counter$count = 6858;
	#10 counter$count = 6859;
	#10 counter$count = 6860;
	#10 counter$count = 6861;
	#10 counter$count = 6862;
	#10 counter$count = 6863;
	#10 counter$count = 6864;
	#10 counter$count = 6865;
	#10 counter$count = 6866;
	#10 counter$count = 6867;
	#10 counter$count = 6868;
	#10 counter$count = 6869;
	#10 counter$count = 6870;
	#10 counter$count = 6871;
	#10 counter$count = 6872;
	#10 counter$count = 6873;
	#10 counter$count = 6874;
	#10 counter$count = 6875;
	#10 counter$count = 6876;
	#10 counter$count = 6877;
	#10 counter$count = 6878;
	#10 counter$count = 6879;
	#10 counter$count = 6880;
	#10 counter$count = 6881;
	#10 counter$count = 6882;
	#10 counter$count = 6883;
	#10 counter$count = 6884;
	#10 counter$count = 6885;
	#10 counter$count = 6886;
	#10 counter$count = 6887;
	#10 counter$count = 6888;
	#10 counter$count = 6889;
	#10 counter$count = 6890;
	#10 counter$count = 6891;
	#10 counter$count = 6892;
	#10 counter$count = 6893;
	#10 counter$count = 6894;
	#10 counter$count = 6895;
	#10 counter$count = 6896;
	#10 counter$count = 6897;
	#10 counter$count = 6898;
	#10 counter$count = 6899;
	#10 counter$count = 6900;
	#10 counter$count = 6901;
	#10 counter$count = 6902;
	#10 counter$count = 6903;
	#10 counter$count = 6904;
	#10 counter$count = 6905;
	#10 counter$count = 6906;
	#10 counter$count = 6907;
	#10 counter$count = 6908;
	#10 counter$count = 6909;
	#10 counter$count = 6910;
	#10 counter$count = 6911;
	#10 counter$count = 6912;
	#10 counter$count = 6913;
	#10 counter$count = 6914;
	#10 counter$count = 6915;
	#10 counter$count = 6916;
	#10 counter$count = 6917;
	#10 counter$count = 6918;
	#10 counter$count = 6919;
	#10 counter$count = 6920;
	#10 counter$count = 6921;
	#10 counter$count = 6922;
	#10 counter$count = 6923;
	#10 counter$count = 6924;
	#10 counter$count = 6925;
	#10 counter$count = 6926;
	#10 counter$count = 6927;
	#10 counter$count = 6928;
	#10 counter$count = 6929;
	#10 counter$count = 6930;
	#10 counter$count = 6931;
	#10 counter$count = 6932;
	#10 counter$count = 6933;
	#10 counter$count = 6934;
	#10 counter$count = 6935;
	#10 counter$count = 6936;
	#10 counter$count = 6937;
	#10 counter$count = 6938;
	#10 counter$count = 6939;
	#10 counter$count = 6940;
	#10 counter$count = 6941;
	#10 counter$count = 6942;
	#10 counter$count = 6943;
	#10 counter$count = 6944;
	#10 counter$count = 6945;
	#10 counter$count = 6946;
	#10 counter$count = 6947;
	#10 counter$count = 6948;
	#10 counter$count = 6949;
	#10 counter$count = 6950;
	#10 counter$count = 6951;
	#10 counter$count = 6952;
	#10 counter$count = 6953;
	#10 counter$count = 6954;
	#10 counter$count = 6955;
	#10 counter$count = 6956;
	#10 counter$count = 6957;
	#10 counter$count = 6958;
	#10 counter$count = 6959;
	#10 counter$count = 6960;
	#10 counter$count = 6961;
	#10 counter$count = 6962;
	#10 counter$count = 6963;
	#10 counter$count = 6964;
	#10 counter$count = 6965;
	#10 counter$count = 6966;
	#10 counter$count = 6967;
	#10 counter$count = 6968;
	#10 counter$count = 6969;
	#10 counter$count = 6970;
	#10 counter$count = 6971;
	#10 counter$count = 6972;
	#10 counter$count = 6973;
	#10 counter$count = 6974;
	#10 counter$count = 6975;
	#10 counter$count = 6976;
	#10 counter$count = 6977;
	#10 counter$count = 6978;
	#10 counter$count = 6979;
	#10 counter$count = 6980;
	#10 counter$count = 6981;
	#10 counter$count = 6982;
	#10 counter$count = 6983;
	#10 counter$count = 6984;
	#10 counter$count = 6985;
	#10 counter$count = 6986;
	#10 counter$count = 6987;
	#10 counter$count = 6988;
	#10 counter$count = 6989;
	#10 counter$count = 6990;
	#10 counter$count = 6991;
	#10 counter$count = 6992;
	#10 counter$count = 6993;
	#10 counter$count = 6994;
	#10 counter$count = 6995;
	#10 counter$count = 6996;
	#10 counter$count = 6997;
	#10 counter$count = 6998;
	#10 counter$count = 6999;
	#10 counter$count = 7000;
	#10 counter$count = 7001;
	#10 counter$count = 7002;
	#10 counter$count = 7003;
	#10 counter$count = 7004;
	#10 counter$count = 7005;
	#10 counter$count = 7006;
	#10 counter$count = 7007;
	#10 counter$count = 7008;
	#10 counter$count = 7009;
	#10 counter$count = 7010;
	#10 counter$count = 7011;
	#10 counter$count = 7012;
	#10 counter$count = 7013;
	#10 counter$count = 7014;
	#10 counter$count = 7015;
	#10 counter$count = 7016;
	#10 counter$count = 7017;
	#10 counter$count = 7018;
	#10 counter$count = 7019;
	#10 counter$count = 7020;
	#10 counter$count = 7021;
	#10 counter$count = 7022;
	#10 counter$count = 7023;
	#10 counter$count = 7024;
	#10 counter$count = 7025;
	#10 counter$count = 7026;
	#10 counter$count = 7027;
	#10 counter$count = 7028;
	#10 counter$count = 7029;
	#10 counter$count = 7030;
	#10 counter$count = 7031;
	#10 counter$count = 7032;
	#10 counter$count = 7033;
	#10 counter$count = 7034;
	#10 counter$count = 7035;
	#10 counter$count = 7036;
	#10 counter$count = 7037;
	#10 counter$count = 7038;
	#10 counter$count = 7039;
	#10 counter$count = 7040;
	#10 counter$count = 7041;
	#10 counter$count = 7042;
	#10 counter$count = 7043;
	#10 counter$count = 7044;
	#10 counter$count = 7045;
	#10 counter$count = 7046;
	#10 counter$count = 7047;
	#10 counter$count = 7048;
	#10 counter$count = 7049;
	#10 counter$count = 7050;
	#10 counter$count = 7051;
	#10 counter$count = 7052;
	#10 counter$count = 7053;
	#10 counter$count = 7054;
	#10 counter$count = 7055;
	#10 counter$count = 7056;
	#10 counter$count = 7057;
	#10 counter$count = 7058;
	#10 counter$count = 7059;
	#10 counter$count = 7060;
	#10 counter$count = 7061;
	#10 counter$count = 7062;
	#10 counter$count = 7063;
	#10 counter$count = 7064;
	#10 counter$count = 7065;
	#10 counter$count = 7066;
	#10 counter$count = 7067;
	#10 counter$count = 7068;
	#10 counter$count = 7069;
	#10 counter$count = 7070;
	#10 counter$count = 7071;
	#10 counter$count = 7072;
	#10 counter$count = 7073;
	#10 counter$count = 7074;
	#10 counter$count = 7075;
	#10 counter$count = 7076;
	#10 counter$count = 7077;
	#10 counter$count = 7078;
	#10 counter$count = 7079;
	#10 counter$count = 7080;
	#10 counter$count = 7081;
	#10 counter$count = 7082;
	#10 counter$count = 7083;
	#10 counter$count = 7084;
	#10 counter$count = 7085;
	#10 counter$count = 7086;
	#10 counter$count = 7087;
	#10 counter$count = 7088;
	#10 counter$count = 7089;
	#10 counter$count = 7090;
	#10 counter$count = 7091;
	#10 counter$count = 7092;
	#10 counter$count = 7093;
	#10 counter$count = 7094;
	#10 counter$count = 7095;
	#10 counter$count = 7096;
	#10 counter$count = 7097;
	#10 counter$count = 7098;
	#10 counter$count = 7099;
	#10 counter$count = 7100;
	#10 counter$count = 7101;
	#10 counter$count = 7102;
	#10 counter$count = 7103;
	#10 counter$count = 7104;
	#10 counter$count = 7105;
	#10 counter$count = 7106;
	#10 counter$count = 7107;
	#10 counter$count = 7108;
	#10 counter$count = 7109;
	#10 counter$count = 7110;
	#10 counter$count = 7111;
	#10 counter$count = 7112;
	#10 counter$count = 7113;
	#10 counter$count = 7114;
	#10 counter$count = 7115;
	#10 counter$count = 7116;
	#10 counter$count = 7117;
	#10 counter$count = 7118;
	#10 counter$count = 7119;
	#10 counter$count = 7120;
	#10 counter$count = 7121;
	#10 counter$count = 7122;
	#10 counter$count = 7123;
	#10 counter$count = 7124;
	#10 counter$count = 7125;
	#10 counter$count = 7126;
	#10 counter$count = 7127;
	#10 counter$count = 7128;
	#10 counter$count = 7129;
	#10 counter$count = 7130;
	#10 counter$count = 7131;
	#10 counter$count = 7132;
	#10 counter$count = 7133;
	#10 counter$count = 7134;
	#10 counter$count = 7135;
	#10 counter$count = 7136;
	#10 counter$count = 7137;
	#10 counter$count = 7138;
	#10 counter$count = 7139;
	#10 counter$count = 7140;
	#10 counter$count = 7141;
	#10 counter$count = 7142;
	#10 counter$count = 7143;
	#10 counter$count = 7144;
	#10 counter$count = 7145;
	#10 counter$count = 7146;
	#10 counter$count = 7147;
	#10 counter$count = 7148;
	#10 counter$count = 7149;
	#10 counter$count = 7150;
	#10 counter$count = 7151;
	#10 counter$count = 7152;
	#10 counter$count = 7153;
	#10 counter$count = 7154;
	#10 counter$count = 7155;
	#10 counter$count = 7156;
	#10 counter$count = 7157;
	#10 counter$count = 7158;
	#10 counter$count = 7159;
	#10 counter$count = 7160;
	#10 counter$count = 7161;
	#10 counter$count = 7162;
	#10 counter$count = 7163;
	#10 counter$count = 7164;
	#10 counter$count = 7165;
	#10 counter$count = 7166;
	#10 counter$count = 7167;
	#10 counter$count = 7168;
	#10 counter$count = 7169;
	#10 counter$count = 7170;
	#10 counter$count = 7171;
	#10 counter$count = 7172;
	#10 counter$count = 7173;
	#10 counter$count = 7174;
	#10 counter$count = 7175;
	#10 counter$count = 7176;
	#10 counter$count = 7177;
	#10 counter$count = 7178;
	#10 counter$count = 7179;
	#10 counter$count = 7180;
	#10 counter$count = 7181;
	#10 counter$count = 7182;
	#10 counter$count = 7183;
	#10 counter$count = 7184;
	#10 counter$count = 7185;
	#10 counter$count = 7186;
	#10 counter$count = 7187;
	#10 counter$count = 7188;
	#10 counter$count = 7189;
	#10 counter$count = 7190;
	#10 counter$count = 7191;
	#10 counter$count = 7192;
	#10 counter$count = 7193;
	#10 counter$count = 7194;
	#10 counter$count = 7195;
	#10 counter$count = 7196;
	#10 counter$count = 7197;
	#10 counter$count = 7198;
	#10 counter$count = 7199;
	#10 counter$count = 7200;
	#10 counter$count = 7201;
	#10 counter$count = 7202;
	#10 counter$count = 7203;
	#10 counter$count = 7204;
	#10 counter$count = 7205;
	#10 counter$count = 7206;
	#10 counter$count = 7207;
	#10 counter$count = 7208;
	#10 counter$count = 7209;
	#10 counter$count = 7210;
	#10 counter$count = 7211;
	#10 counter$count = 7212;
	#10 counter$count = 7213;
	#10 counter$count = 7214;
	#10 counter$count = 7215;
	#10 counter$count = 7216;
	#10 counter$count = 7217;
	#10 counter$count = 7218;
	#10 counter$count = 7219;
	#10 counter$count = 7220;
	#10 counter$count = 7221;
	#10 counter$count = 7222;
	#10 counter$count = 7223;
	#10 counter$count = 7224;
	#10 counter$count = 7225;
	#10 counter$count = 7226;
	#10 counter$count = 7227;
	#10 counter$count = 7228;
	#10 counter$count = 7229;
	#10 counter$count = 7230;
	#10 counter$count = 7231;
	#10 counter$count = 7232;
	#10 counter$count = 7233;
	#10 counter$count = 7234;
	#10 counter$count = 7235;
	#10 counter$count = 7236;
	#10 counter$count = 7237;
	#10 counter$count = 7238;
	#10 counter$count = 7239;
	#10 counter$count = 7240;
	#10 counter$count = 7241;
	#10 counter$count = 7242;
	#10 counter$count = 7243;
	#10 counter$count = 7244;
	#10 counter$count = 7245;
	#10 counter$count = 7246;
	#10 counter$count = 7247;
	#10 counter$count = 7248;
	#10 counter$count = 7249;
	#10 counter$count = 7250;
	#10 counter$count = 7251;
	#10 counter$count = 7252;
	#10 counter$count = 7253;
	#10 counter$count = 7254;
	#10 counter$count = 7255;
	#10 counter$count = 7256;
	#10 counter$count = 7257;
	#10 counter$count = 7258;
	#10 counter$count = 7259;
	#10 counter$count = 7260;
	#10 counter$count = 7261;
	#10 counter$count = 7262;
	#10 counter$count = 7263;
	#10 counter$count = 7264;
	#10 counter$count = 7265;
	#10 counter$count = 7266;
	#10 counter$count = 7267;
	#10 counter$count = 7268;
	#10 counter$count = 7269;
	#10 counter$count = 7270;
	#10 counter$count = 7271;
	#10 counter$count = 7272;
	#10 counter$count = 7273;
	#10 counter$count = 7274;
	#10 counter$count = 7275;
	#10 counter$count = 7276;
	#10 counter$count = 7277;
	#10 counter$count = 7278;
	#10 counter$count = 7279;
	#10 counter$count = 7280;
	#10 counter$count = 7281;
	#10 counter$count = 7282;
	#10 counter$count = 7283;
	#10 counter$count = 7284;
	#10 counter$count = 7285;
	#10 counter$count = 7286;
	#10 counter$count = 7287;
	#10 counter$count = 7288;
	#10 counter$count = 7289;
	#10 counter$count = 7290;
	#10 counter$count = 7291;
	#10 counter$count = 7292;
	#10 counter$count = 7293;
	#10 counter$count = 7294;
	#10 counter$count = 7295;
	#10 counter$count = 7296;
	#10 counter$count = 7297;
	#10 counter$count = 7298;
	#10 counter$count = 7299;
	#10 counter$count = 7300;
	#10 counter$count = 7301;
	#10 counter$count = 7302;
	#10 counter$count = 7303;
	#10 counter$count = 7304;
	#10 counter$count = 7305;
	#10 counter$count = 7306;
	#10 counter$count = 7307;
	#10 counter$count = 7308;
	#10 counter$count = 7309;
	#10 counter$count = 7310;
	#10 counter$count = 7311;
	#10 counter$count = 7312;
	#10 counter$count = 7313;
	#10 counter$count = 7314;
	#10 counter$count = 7315;
	#10 counter$count = 7316;
	#10 counter$count = 7317;
	#10 counter$count = 7318;
	#10 counter$count = 7319;
	#10 counter$count = 7320;
	#10 counter$count = 7321;
	#10 counter$count = 7322;
	#10 counter$count = 7323;
	#10 counter$count = 7324;
	#10 counter$count = 7325;
	#10 counter$count = 7326;
	#10 counter$count = 7327;
	#10 counter$count = 7328;
	#10 counter$count = 7329;
	#10 counter$count = 7330;
	#10 counter$count = 7331;
	#10 counter$count = 7332;
	#10 counter$count = 7333;
	#10 counter$count = 7334;
	#10 counter$count = 7335;
	#10 counter$count = 7336;
	#10 counter$count = 7337;
	#10 counter$count = 7338;
	#10 counter$count = 7339;
	#10 counter$count = 7340;
	#10 counter$count = 7341;
	#10 counter$count = 7342;
	#10 counter$count = 7343;
	#10 counter$count = 7344;
	#10 counter$count = 7345;
	#10 counter$count = 7346;
	#10 counter$count = 7347;
	#10 counter$count = 7348;
	#10 counter$count = 7349;
	#10 counter$count = 7350;
	#10 counter$count = 7351;
	#10 counter$count = 7352;
	#10 counter$count = 7353;
	#10 counter$count = 7354;
	#10 counter$count = 7355;
	#10 counter$count = 7356;
	#10 counter$count = 7357;
	#10 counter$count = 7358;
	#10 counter$count = 7359;
	#10 counter$count = 7360;
	#10 counter$count = 7361;
	#10 counter$count = 7362;
	#10 counter$count = 7363;
	#10 counter$count = 7364;
	#10 counter$count = 7365;
	#10 counter$count = 7366;
	#10 counter$count = 7367;
	#10 counter$count = 7368;
	#10 counter$count = 7369;
	#10 counter$count = 7370;
	#10 counter$count = 7371;
	#10 counter$count = 7372;
	#10 counter$count = 7373;
	#10 counter$count = 7374;
	#10 counter$count = 7375;
	#10 counter$count = 7376;
	#10 counter$count = 7377;
	#10 counter$count = 7378;
	#10 counter$count = 7379;
	#10 counter$count = 7380;
	#10 counter$count = 7381;
	#10 counter$count = 7382;
	#10 counter$count = 7383;
	#10 counter$count = 7384;
	#10 counter$count = 7385;
	#10 counter$count = 7386;
	#10 counter$count = 7387;
	#10 counter$count = 7388;
	#10 counter$count = 7389;
	#10 counter$count = 7390;
	#10 counter$count = 7391;
	#10 counter$count = 7392;
	#10 counter$count = 7393;
	#10 counter$count = 7394;
	#10 counter$count = 7395;
	#10 counter$count = 7396;
	#10 counter$count = 7397;
	#10 counter$count = 7398;
	#10 counter$count = 7399;
	#10 counter$count = 7400;
	#10 counter$count = 7401;
	#10 counter$count = 7402;
	#10 counter$count = 7403;
	#10 counter$count = 7404;
	#10 counter$count = 7405;
	#10 counter$count = 7406;
	#10 counter$count = 7407;
	#10 counter$count = 7408;
	#10 counter$count = 7409;
	#10 counter$count = 7410;
	#10 counter$count = 7411;
	#10 counter$count = 7412;
	#10 counter$count = 7413;
	#10 counter$count = 7414;
	#10 counter$count = 7415;
	#10 counter$count = 7416;
	#10 counter$count = 7417;
	#10 counter$count = 7418;
	#10 counter$count = 7419;
	#10 counter$count = 7420;
	#10 counter$count = 7421;
	#10 counter$count = 7422;
	#10 counter$count = 7423;
	#10 counter$count = 7424;
	#10 counter$count = 7425;
	#10 counter$count = 7426;
	#10 counter$count = 7427;
	#10 counter$count = 7428;
	#10 counter$count = 7429;
	#10 counter$count = 7430;
	#10 counter$count = 7431;
	#10 counter$count = 7432;
	#10 counter$count = 7433;
	#10 counter$count = 7434;
	#10 counter$count = 7435;
	#10 counter$count = 7436;
	#10 counter$count = 7437;
	#10 counter$count = 7438;
	#10 counter$count = 7439;
	#10 counter$count = 7440;
	#10 counter$count = 7441;
	#10 counter$count = 7442;
	#10 counter$count = 7443;
	#10 counter$count = 7444;
	#10 counter$count = 7445;
	#10 counter$count = 7446;
	#10 counter$count = 7447;
	#10 counter$count = 7448;
	#10 counter$count = 7449;
	#10 counter$count = 7450;
	#10 counter$count = 7451;
	#10 counter$count = 7452;
	#10 counter$count = 7453;
	#10 counter$count = 7454;
	#10 counter$count = 7455;
	#10 counter$count = 7456;
	#10 counter$count = 7457;
	#10 counter$count = 7458;
	#10 counter$count = 7459;
	#10 counter$count = 7460;
	#10 counter$count = 7461;
	#10 counter$count = 7462;
	#10 counter$count = 7463;
	#10 counter$count = 7464;
	#10 counter$count = 7465;
	#10 counter$count = 7466;
	#10 counter$count = 7467;
	#10 counter$count = 7468;
	#10 counter$count = 7469;
	#10 counter$count = 7470;
	#10 counter$count = 7471;
	#10 counter$count = 7472;
	#10 counter$count = 7473;
	#10 counter$count = 7474;
	#10 counter$count = 7475;
	#10 counter$count = 7476;
	#10 counter$count = 7477;
	#10 counter$count = 7478;
	#10 counter$count = 7479;
	#10 counter$count = 7480;
	#10 counter$count = 7481;
	#10 counter$count = 7482;
	#10 counter$count = 7483;
	#10 counter$count = 7484;
	#10 counter$count = 7485;
	#10 counter$count = 7486;
	#10 counter$count = 7487;
	#10 counter$count = 7488;
	#10 counter$count = 7489;
	#10 counter$count = 7490;
	#10 counter$count = 7491;
	#10 counter$count = 7492;
	#10 counter$count = 7493;
	#10 counter$count = 7494;
	#10 counter$count = 7495;
	#10 counter$count = 7496;
	#10 counter$count = 7497;
	#10 counter$count = 7498;
	#10 counter$count = 7499;
	#10 counter$count = 7500;
	#10 counter$count = 7501;
	#10 counter$count = 7502;
	#10 counter$count = 7503;
	#10 counter$count = 7504;
	#10 counter$count = 7505;
	#10 counter$count = 7506;
	#10 counter$count = 7507;
	#10 counter$count = 7508;
	#10 counter$count = 7509;
	#10 counter$count = 7510;
	#10 counter$count = 7511;
	#10 counter$count = 7512;
	#10 counter$count = 7513;
	#10 counter$count = 7514;
	#10 counter$count = 7515;
	#10 counter$count = 7516;
	#10 counter$count = 7517;
	#10 counter$count = 7518;
	#10 counter$count = 7519;
	#10 counter$count = 7520;
	#10 counter$count = 7521;
	#10 counter$count = 7522;
	#10 counter$count = 7523;
	#10 counter$count = 7524;
	#10 counter$count = 7525;
	#10 counter$count = 7526;
	#10 counter$count = 7527;
	#10 counter$count = 7528;
	#10 counter$count = 7529;
	#10 counter$count = 7530;
	#10 counter$count = 7531;
	#10 counter$count = 7532;
	#10 counter$count = 7533;
	#10 counter$count = 7534;
	#10 counter$count = 7535;
	#10 counter$count = 7536;
	#10 counter$count = 7537;
	#10 counter$count = 7538;
	#10 counter$count = 7539;
	#10 counter$count = 7540;
	#10 counter$count = 7541;
	#10 counter$count = 7542;
	#10 counter$count = 7543;
	#10 counter$count = 7544;
	#10 counter$count = 7545;
	#10 counter$count = 7546;
	#10 counter$count = 7547;
	#10 counter$count = 7548;
	#10 counter$count = 7549;
	#10 counter$count = 7550;
	#10 counter$count = 7551;
	#10 counter$count = 7552;
	#10 counter$count = 7553;
	#10 counter$count = 7554;
	#10 counter$count = 7555;
	#10 counter$count = 7556;
	#10 counter$count = 7557;
	#10 counter$count = 7558;
	#10 counter$count = 7559;
	#10 counter$count = 7560;
	#10 counter$count = 7561;
	#10 counter$count = 7562;
	#10 counter$count = 7563;
	#10 counter$count = 7564;
	#10 counter$count = 7565;
	#10 counter$count = 7566;
	#10 counter$count = 7567;
	#10 counter$count = 7568;
	#10 counter$count = 7569;
	#10 counter$count = 7570;
	#10 counter$count = 7571;
	#10 counter$count = 7572;
	#10 counter$count = 7573;
	#10 counter$count = 7574;
	#10 counter$count = 7575;
	#10 counter$count = 7576;
	#10 counter$count = 7577;
	#10 counter$count = 7578;
	#10 counter$count = 7579;
	#10 counter$count = 7580;
	#10 counter$count = 7581;
	#10 counter$count = 7582;
	#10 counter$count = 7583;
	#10 counter$count = 7584;
	#10 counter$count = 7585;
	#10 counter$count = 7586;
	#10 counter$count = 7587;
	#10 counter$count = 7588;
	#10 counter$count = 7589;
	#10 counter$count = 7590;
	#10 counter$count = 7591;
	#10 counter$count = 7592;
	#10 counter$count = 7593;
	#10 counter$count = 7594;
	#10 counter$count = 7595;
	#10 counter$count = 7596;
	#10 counter$count = 7597;
	#10 counter$count = 7598;
	#10 counter$count = 7599;
	#10 counter$count = 7600;
	#10 counter$count = 7601;
	#10 counter$count = 7602;
	#10 counter$count = 7603;
	#10 counter$count = 7604;
	#10 counter$count = 7605;
	#10 counter$count = 7606;
	#10 counter$count = 7607;
	#10 counter$count = 7608;
	#10 counter$count = 7609;
	#10 counter$count = 7610;
	#10 counter$count = 7611;
	#10 counter$count = 7612;
	#10 counter$count = 7613;
	#10 counter$count = 7614;
	#10 counter$count = 7615;
	#10 counter$count = 7616;
	#10 counter$count = 7617;
	#10 counter$count = 7618;
	#10 counter$count = 7619;
	#10 counter$count = 7620;
	#10 counter$count = 7621;
	#10 counter$count = 7622;
	#10 counter$count = 7623;
	#10 counter$count = 7624;
	#10 counter$count = 7625;
	#10 counter$count = 7626;
	#10 counter$count = 7627;
	#10 counter$count = 7628;
	#10 counter$count = 7629;
	#10 counter$count = 7630;
	#10 counter$count = 7631;
	#10 counter$count = 7632;
	#10 counter$count = 7633;
	#10 counter$count = 7634;
	#10 counter$count = 7635;
	#10 counter$count = 7636;
	#10 counter$count = 7637;
	#10 counter$count = 7638;
	#10 counter$count = 7639;
	#10 counter$count = 7640;
	#10 counter$count = 7641;
	#10 counter$count = 7642;
	#10 counter$count = 7643;
	#10 counter$count = 7644;
	#10 counter$count = 7645;
	#10 counter$count = 7646;
	#10 counter$count = 7647;
	#10 counter$count = 7648;
	#10 counter$count = 7649;
	#10 counter$count = 7650;
	#10 counter$count = 7651;
	#10 counter$count = 7652;
	#10 counter$count = 7653;
	#10 counter$count = 7654;
	#10 counter$count = 7655;
	#10 counter$count = 7656;
	#10 counter$count = 7657;
	#10 counter$count = 7658;
	#10 counter$count = 7659;
	#10 counter$count = 7660;
	#10 counter$count = 7661;
	#10 counter$count = 7662;
	#10 counter$count = 7663;
	#10 counter$count = 7664;
	#10 counter$count = 7665;
	#10 counter$count = 7666;
	#10 counter$count = 7667;
	#10 counter$count = 7668;
	#10 counter$count = 7669;
	#10 counter$count = 7670;
	#10 counter$count = 7671;
	#10 counter$count = 7672;
	#10 counter$count = 7673;
	#10 counter$count = 7674;
	#10 counter$count = 7675;
	#10 counter$count = 7676;
	#10 counter$count = 7677;
	#10 counter$count = 7678;
	#10 counter$count = 7679;
	#10 counter$count = 7680;
	#10 counter$count = 7681;
	#10 counter$count = 7682;
	#10 counter$count = 7683;
	#10 counter$count = 7684;
	#10 counter$count = 7685;
	#10 counter$count = 7686;
	#10 counter$count = 7687;
	#10 counter$count = 7688;
	#10 counter$count = 7689;
	#10 counter$count = 7690;
	#10 counter$count = 7691;
	#10 counter$count = 7692;
	#10 counter$count = 7693;
	#10 counter$count = 7694;
	#10 counter$count = 7695;
	#10 counter$count = 7696;
	#10 counter$count = 7697;
	#10 counter$count = 7698;
	#10 counter$count = 7699;
	#10 counter$count = 7700;
	#10 counter$count = 7701;
	#10 counter$count = 7702;
	#10 counter$count = 7703;
	#10 counter$count = 7704;
	#10 counter$count = 7705;
	#10 counter$count = 7706;
	#10 counter$count = 7707;
	#10 counter$count = 7708;
	#10 counter$count = 7709;
	#10 counter$count = 7710;
	#10 counter$count = 7711;
	#10 counter$count = 7712;
	#10 counter$count = 7713;
	#10 counter$count = 7714;
	#10 counter$count = 7715;
	#10 counter$count = 7716;
	#10 counter$count = 7717;
	#10 counter$count = 7718;
	#10 counter$count = 7719;
	#10 counter$count = 7720;
	#10 counter$count = 7721;
	#10 counter$count = 7722;
	#10 counter$count = 7723;
	#10 counter$count = 7724;
	#10 counter$count = 7725;
	#10 counter$count = 7726;
	#10 counter$count = 7727;
	#10 counter$count = 7728;
	#10 counter$count = 7729;
	#10 counter$count = 7730;
	#10 counter$count = 7731;
	#10 counter$count = 7732;
	#10 counter$count = 7733;
	#10 counter$count = 7734;
	#10 counter$count = 7735;
	#10 counter$count = 7736;
	#10 counter$count = 7737;
	#10 counter$count = 7738;
	#10 counter$count = 7739;
	#10 counter$count = 7740;
	#10 counter$count = 7741;
	#10 counter$count = 7742;
	#10 counter$count = 7743;
	#10 counter$count = 7744;
	#10 counter$count = 7745;
	#10 counter$count = 7746;
	#10 counter$count = 7747;
	#10 counter$count = 7748;
	#10 counter$count = 7749;
	#10 counter$count = 7750;
	#10 counter$count = 7751;
	#10 counter$count = 7752;
	#10 counter$count = 7753;
	#10 counter$count = 7754;
	#10 counter$count = 7755;
	#10 counter$count = 7756;
	#10 counter$count = 7757;
	#10 counter$count = 7758;
	#10 counter$count = 7759;
	#10 counter$count = 7760;
	#10 counter$count = 7761;
	#10 counter$count = 7762;
	#10 counter$count = 7763;
	#10 counter$count = 7764;
	#10 counter$count = 7765;
	#10 counter$count = 7766;
	#10 counter$count = 7767;
	#10 counter$count = 7768;
	#10 counter$count = 7769;
	#10 counter$count = 7770;
	#10 counter$count = 7771;
	#10 counter$count = 7772;
	#10 counter$count = 7773;
	#10 counter$count = 7774;
	#10 counter$count = 7775;
	#10 counter$count = 7776;
	#10 counter$count = 7777;
	#10 counter$count = 7778;
	#10 counter$count = 7779;
	#10 counter$count = 7780;
	#10 counter$count = 7781;
	#10 counter$count = 7782;
	#10 counter$count = 7783;
	#10 counter$count = 7784;
	#10 counter$count = 7785;
	#10 counter$count = 7786;
	#10 counter$count = 7787;
	#10 counter$count = 7788;
	#10 counter$count = 7789;
	#10 counter$count = 7790;
	#10 counter$count = 7791;
	#10 counter$count = 7792;
	#10 counter$count = 7793;
	#10 counter$count = 7794;
	#10 counter$count = 7795;
	#10 counter$count = 7796;
	#10 counter$count = 7797;
	#10 counter$count = 7798;
	#10 counter$count = 7799;
	#10 counter$count = 7800;
	#10 counter$count = 7801;
	#10 counter$count = 7802;
	#10 counter$count = 7803;
	#10 counter$count = 7804;
	#10 counter$count = 7805;
	#10 counter$count = 7806;
	#10 counter$count = 7807;
	#10 counter$count = 7808;
	#10 counter$count = 7809;
	#10 counter$count = 7810;
	#10 counter$count = 7811;
	#10 counter$count = 7812;
	#10 counter$count = 7813;
	#10 counter$count = 7814;
	#10 counter$count = 7815;
	#10 counter$count = 7816;
	#10 counter$count = 7817;
	#10 counter$count = 7818;
	#10 counter$count = 7819;
	#10 counter$count = 7820;
	#10 counter$count = 7821;
	#10 counter$count = 7822;
	#10 counter$count = 7823;
	#10 counter$count = 7824;
	#10 counter$count = 7825;
	#10 counter$count = 7826;
	#10 counter$count = 7827;
	#10 counter$count = 7828;
	#10 counter$count = 7829;
	#10 counter$count = 7830;
	#10 counter$count = 7831;
	#10 counter$count = 7832;
	#10 counter$count = 7833;
	#10 counter$count = 7834;
	#10 counter$count = 7835;
	#10 counter$count = 7836;
	#10 counter$count = 7837;
	#10 counter$count = 7838;
	#10 counter$count = 7839;
	#10 counter$count = 7840;
	#10 counter$count = 7841;
	#10 counter$count = 7842;
	#10 counter$count = 7843;
	#10 counter$count = 7844;
	#10 counter$count = 7845;
	#10 counter$count = 7846;
	#10 counter$count = 7847;
	#10 counter$count = 7848;
	#10 counter$count = 7849;
	#10 counter$count = 7850;
	#10 counter$count = 7851;
	#10 counter$count = 7852;
	#10 counter$count = 7853;
	#10 counter$count = 7854;
	#10 counter$count = 7855;
	#10 counter$count = 7856;
	#10 counter$count = 7857;
	#10 counter$count = 7858;
	#10 counter$count = 7859;
	#10 counter$count = 7860;
	#10 counter$count = 7861;
	#10 counter$count = 7862;
	#10 counter$count = 7863;
	#10 counter$count = 7864;
	#10 counter$count = 7865;
	#10 counter$count = 7866;
	#10 counter$count = 7867;
	#10 counter$count = 7868;
	#10 counter$count = 7869;
	#10 counter$count = 7870;
	#10 counter$count = 7871;
	#10 counter$count = 7872;
	#10 counter$count = 7873;
	#10 counter$count = 7874;
	#10 counter$count = 7875;
	#10 counter$count = 7876;
	#10 counter$count = 7877;
	#10 counter$count = 7878;
	#10 counter$count = 7879;
	#10 counter$count = 7880;
	#10 counter$count = 7881;
	#10 counter$count = 7882;
	#10 counter$count = 7883;
	#10 counter$count = 7884;
	#10 counter$count = 7885;
	#10 counter$count = 7886;
	#10 counter$count = 7887;
	#10 counter$count = 7888;
	#10 counter$count = 7889;
	#10 counter$count = 7890;
	#10 counter$count = 7891;
	#10 counter$count = 7892;
	#10 counter$count = 7893;
	#10 counter$count = 7894;
	#10 counter$count = 7895;
	#10 counter$count = 7896;
	#10 counter$count = 7897;
	#10 counter$count = 7898;
	#10 counter$count = 7899;
	#10 counter$count = 7900;
	#10 counter$count = 7901;
	#10 counter$count = 7902;
	#10 counter$count = 7903;
	#10 counter$count = 7904;
	#10 counter$count = 7905;
	#10 counter$count = 7906;
	#10 counter$count = 7907;
	#10 counter$count = 7908;
	#10 counter$count = 7909;
	#10 counter$count = 7910;
	#10 counter$count = 7911;
	#10 counter$count = 7912;
	#10 counter$count = 7913;
	#10 counter$count = 7914;
	#10 counter$count = 7915;
	#10 counter$count = 7916;
	#10 counter$count = 7917;
	#10 counter$count = 7918;
	#10 counter$count = 7919;
	#10 counter$count = 7920;
	#10 counter$count = 7921;
	#10 counter$count = 7922;
	#10 counter$count = 7923;
	#10 counter$count = 7924;
	#10 counter$count = 7925;
	#10 counter$count = 7926;
	#10 counter$count = 7927;
	#10 counter$count = 7928;
	#10 counter$count = 7929;
	#10 counter$count = 7930;
	#10 counter$count = 7931;
	#10 counter$count = 7932;
	#10 counter$count = 7933;
	#10 counter$count = 7934;
	#10 counter$count = 7935;
	#10 counter$count = 7936;
	#10 counter$count = 7937;
	#10 counter$count = 7938;
	#10 counter$count = 7939;
	#10 counter$count = 7940;
	#10 counter$count = 7941;
	#10 counter$count = 7942;
	#10 counter$count = 7943;
	#10 counter$count = 7944;
	#10 counter$count = 7945;
	#10 counter$count = 7946;
	#10 counter$count = 7947;
	#10 counter$count = 7948;
	#10 counter$count = 7949;
	#10 counter$count = 7950;
	#10 counter$count = 7951;
	#10 counter$count = 7952;
	#10 counter$count = 7953;
	#10 counter$count = 7954;
	#10 counter$count = 7955;
	#10 counter$count = 7956;
	#10 counter$count = 7957;
	#10 counter$count = 7958;
	#10 counter$count = 7959;
	#10 counter$count = 7960;
	#10 counter$count = 7961;
	#10 counter$count = 7962;
	#10 counter$count = 7963;
	#10 counter$count = 7964;
	#10 counter$count = 7965;
	#10 counter$count = 7966;
	#10 counter$count = 7967;
	#10 counter$count = 7968;
	#10 counter$count = 7969;
	#10 counter$count = 7970;
	#10 counter$count = 7971;
	#10 counter$count = 7972;
	#10 counter$count = 7973;
	#10 counter$count = 7974;
	#10 counter$count = 7975;
	#10 counter$count = 7976;
	#10 counter$count = 7977;
	#10 counter$count = 7978;
	#10 counter$count = 7979;
	#10 counter$count = 7980;
	#10 counter$count = 7981;
	#10 counter$count = 7982;
	#10 counter$count = 7983;
	#10 counter$count = 7984;
	#10 counter$count = 7985;
	#10 counter$count = 7986;
	#10 counter$count = 7987;
	#10 counter$count = 7988;
	#10 counter$count = 7989;
	#10 counter$count = 7990;
	#10 counter$count = 7991;
	#10 counter$count = 7992;
	#10 counter$count = 7993;
	#10 counter$count = 7994;
	#10 counter$count = 7995;
	#10 counter$count = 7996;
	#10 counter$count = 7997;
	#10 counter$count = 7998;
	#10 counter$count = 7999;
	#10 counter$count = 8000;
	#10 counter$count = 8001;
	#10 counter$count = 8002;
	#10 counter$count = 8003;
	#10 counter$count = 8004;
	#10 counter$count = 8005;
	#10 counter$count = 8006;
	#10 counter$count = 8007;
	#10 counter$count = 8008;
	#10 counter$count = 8009;
	#10 counter$count = 8010;
	#10 counter$count = 8011;
	#10 counter$count = 8012;
	#10 counter$count = 8013;
	#10 counter$count = 8014;
	#10 counter$count = 8015;
	#10 counter$count = 8016;
	#10 counter$count = 8017;
	#10 counter$count = 8018;
	#10 counter$count = 8019;
	#10 counter$count = 8020;
	#10 counter$count = 8021;
	#10 counter$count = 8022;
	#10 counter$count = 8023;
	#10 counter$count = 8024;
	#10 counter$count = 8025;
	#10 counter$count = 8026;
	#10 counter$count = 8027;
	#10 counter$count = 8028;
	#10 counter$count = 8029;
	#10 counter$count = 8030;
	#10 counter$count = 8031;
	#10 counter$count = 8032;
	#10 counter$count = 8033;
	#10 counter$count = 8034;
	#10 counter$count = 8035;
	#10 counter$count = 8036;
	#10 counter$count = 8037;
	#10 counter$count = 8038;
	#10 counter$count = 8039;
	#10 counter$count = 8040;
	#10 counter$count = 8041;
	#10 counter$count = 8042;
	#10 counter$count = 8043;
	#10 counter$count = 8044;
	#10 counter$count = 8045;
	#10 counter$count = 8046;
	#10 counter$count = 8047;
	#10 counter$count = 8048;
	#10 counter$count = 8049;
	#10 counter$count = 8050;
	#10 counter$count = 8051;
	#10 counter$count = 8052;
	#10 counter$count = 8053;
	#10 counter$count = 8054;
	#10 counter$count = 8055;
	#10 counter$count = 8056;
	#10 counter$count = 8057;
	#10 counter$count = 8058;
	#10 counter$count = 8059;
	#10 counter$count = 8060;
	#10 counter$count = 8061;
	#10 counter$count = 8062;
	#10 counter$count = 8063;
	#10 counter$count = 8064;
	#10 counter$count = 8065;
	#10 counter$count = 8066;
	#10 counter$count = 8067;
	#10 counter$count = 8068;
	#10 counter$count = 8069;
	#10 counter$count = 8070;
	#10 counter$count = 8071;
	#10 counter$count = 8072;
	#10 counter$count = 8073;
	#10 counter$count = 8074;
	#10 counter$count = 8075;
	#10 counter$count = 8076;
	#10 counter$count = 8077;
	#10 counter$count = 8078;
	#10 counter$count = 8079;
	#10 counter$count = 8080;
	#10 counter$count = 8081;
	#10 counter$count = 8082;
	#10 counter$count = 8083;
	#10 counter$count = 8084;
	#10 counter$count = 8085;
	#10 counter$count = 8086;
	#10 counter$count = 8087;
	#10 counter$count = 8088;
	#10 counter$count = 8089;
	#10 counter$count = 8090;
	#10 counter$count = 8091;
	#10 counter$count = 8092;
	#10 counter$count = 8093;
	#10 counter$count = 8094;
	#10 counter$count = 8095;
	#10 counter$count = 8096;
	#10 counter$count = 8097;
	#10 counter$count = 8098;
	#10 counter$count = 8099;
	#10 counter$count = 8100;
	#10 counter$count = 8101;
	#10 counter$count = 8102;
	#10 counter$count = 8103;
	#10 counter$count = 8104;
	#10 counter$count = 8105;
	#10 counter$count = 8106;
	#10 counter$count = 8107;
	#10 counter$count = 8108;
	#10 counter$count = 8109;
	#10 counter$count = 8110;
	#10 counter$count = 8111;
	#10 counter$count = 8112;
	#10 counter$count = 8113;
	#10 counter$count = 8114;
	#10 counter$count = 8115;
	#10 counter$count = 8116;
	#10 counter$count = 8117;
	#10 counter$count = 8118;
	#10 counter$count = 8119;
	#10 counter$count = 8120;
	#10 counter$count = 8121;
	#10 counter$count = 8122;
	#10 counter$count = 8123;
	#10 counter$count = 8124;
	#10 counter$count = 8125;
	#10 counter$count = 8126;
	#10 counter$count = 8127;
	#10 counter$count = 8128;
	#10 counter$count = 8129;
	#10 counter$count = 8130;
	#10 counter$count = 8131;
	#10 counter$count = 8132;
	#10 counter$count = 8133;
	#10 counter$count = 8134;
	#10 counter$count = 8135;
	#10 counter$count = 8136;
	#10 counter$count = 8137;
	#10 counter$count = 8138;
	#10 counter$count = 8139;
	#10 counter$count = 8140;
	#10 counter$count = 8141;
	#10 counter$count = 8142;
	#10 counter$count = 8143;
	#10 counter$count = 8144;
	#10 counter$count = 8145;
	#10 counter$count = 8146;
	#10 counter$count = 8147;
	#10 counter$count = 8148;
	#10 counter$count = 8149;
	#10 counter$count = 8150;
	#10 counter$count = 8151;
	#10 counter$count = 8152;
	#10 counter$count = 8153;
	#10 counter$count = 8154;
	#10 counter$count = 8155;
	#10 counter$count = 8156;
	#10 counter$count = 8157;
	#10 counter$count = 8158;
	#10 counter$count = 8159;
	#10 counter$count = 8160;
	#10 counter$count = 8161;
	#10 counter$count = 8162;
	#10 counter$count = 8163;
	#10 counter$count = 8164;
	#10 counter$count = 8165;
	#10 counter$count = 8166;
	#10 counter$count = 8167;
	#10 counter$count = 8168;
	#10 counter$count = 8169;
	#10 counter$count = 8170;
	#10 counter$count = 8171;
	#10 counter$count = 8172;
	#10 counter$count = 8173;
	#10 counter$count = 8174;
	#10 counter$count = 8175;
	#10 counter$count = 8176;
	#10 counter$count = 8177;
	#10 counter$count = 8178;
	#10 counter$count = 8179;
	#10 counter$count = 8180;
	#10 counter$count = 8181;
	#10 counter$count = 8182;
	#10 counter$count = 8183;
	#10 counter$count = 8184;
	#10 counter$count = 8185;
	#10 counter$count = 8186;
	#10 counter$count = 8187;
	#10 counter$count = 8188;
	#10 counter$count = 8189;
	#10 counter$count = 8190;
	#10 counter$count = 8191;
	#10 counter$count = 8192;
	#10 counter$count = 8193;
	#10 counter$count = 8194;
	#10 counter$count = 8195;
	#10 counter$count = 8196;
	#10 counter$count = 8197;
	#10 counter$count = 8198;
	#10 counter$count = 8199;
	#10 counter$count = 8200;
	#10 counter$count = 8201;
	#10 counter$count = 8202;
	#10 counter$count = 8203;
	#10 counter$count = 8204;
	#10 counter$count = 8205;
	#10 counter$count = 8206;
	#10 counter$count = 8207;
	#10 counter$count = 8208;
	#10 counter$count = 8209;
	#10 counter$count = 8210;
	#10 counter$count = 8211;
	#10 counter$count = 8212;
	#10 counter$count = 8213;
	#10 counter$count = 8214;
	#10 counter$count = 8215;
	#10 counter$count = 8216;
	#10 counter$count = 8217;
	#10 counter$count = 8218;
	#10 counter$count = 8219;
	#10 counter$count = 8220;
	#10 counter$count = 8221;
	#10 counter$count = 8222;
	#10 counter$count = 8223;
	#10 counter$count = 8224;
	#10 counter$count = 8225;
	#10 counter$count = 8226;
	#10 counter$count = 8227;
	#10 counter$count = 8228;
	#10 counter$count = 8229;
	#10 counter$count = 8230;
	#10 counter$count = 8231;
	#10 counter$count = 8232;
	#10 counter$count = 8233;
	#10 counter$count = 8234;
	#10 counter$count = 8235;
	#10 counter$count = 8236;
	#10 counter$count = 8237;
	#10 counter$count = 8238;
	#10 counter$count = 8239;
	#10 counter$count = 8240;
	#10 counter$count = 8241;
	#10 counter$count = 8242;
	#10 counter$count = 8243;
	#10 counter$count = 8244;
	#10 counter$count = 8245;
	#10 counter$count = 8246;
	#10 counter$count = 8247;
	#10 counter$count = 8248;
	#10 counter$count = 8249;
	#10 counter$count = 8250;
	#10 counter$count = 8251;
	#10 counter$count = 8252;
	#10 counter$count = 8253;
	#10 counter$count = 8254;
	#10 counter$count = 8255;
	#10 counter$count = 8256;
	#10 counter$count = 8257;
	#10 counter$count = 8258;
	#10 counter$count = 8259;
	#10 counter$count = 8260;
	#10 counter$count = 8261;
	#10 counter$count = 8262;
	#10 counter$count = 8263;
	#10 counter$count = 8264;
	#10 counter$count = 8265;
	#10 counter$count = 8266;
	#10 counter$count = 8267;
	#10 counter$count = 8268;
	#10 counter$count = 8269;
	#10 counter$count = 8270;
	#10 counter$count = 8271;
	#10 counter$count = 8272;
	#10 counter$count = 8273;
	#10 counter$count = 8274;
	#10 counter$count = 8275;
	#10 counter$count = 8276;
	#10 counter$count = 8277;
	#10 counter$count = 8278;
	#10 counter$count = 8279;
	#10 counter$count = 8280;
	#10 counter$count = 8281;
	#10 counter$count = 8282;
	#10 counter$count = 8283;
	#10 counter$count = 8284;
	#10 counter$count = 8285;
	#10 counter$count = 8286;
	#10 counter$count = 8287;
	#10 counter$count = 8288;
	#10 counter$count = 8289;
	#10 counter$count = 8290;
	#10 counter$count = 8291;
	#10 counter$count = 8292;
	#10 counter$count = 8293;
	#10 counter$count = 8294;
	#10 counter$count = 8295;
	#10 counter$count = 8296;
	#10 counter$count = 8297;
	#10 counter$count = 8298;
	#10 counter$count = 8299;
	#10 counter$count = 8300;
	#10 counter$count = 8301;
	#10 counter$count = 8302;
	#10 counter$count = 8303;
	#10 counter$count = 8304;
	#10 counter$count = 8305;
	#10 counter$count = 8306;
	#10 counter$count = 8307;
	#10 counter$count = 8308;
	#10 counter$count = 8309;
	#10 counter$count = 8310;
	#10 counter$count = 8311;
	#10 counter$count = 8312;
	#10 counter$count = 8313;
	#10 counter$count = 8314;
	#10 counter$count = 8315;
	#10 counter$count = 8316;
	#10 counter$count = 8317;
	#10 counter$count = 8318;
	#10 counter$count = 8319;
	#10 counter$count = 8320;
	#10 counter$count = 8321;
	#10 counter$count = 8322;
	#10 counter$count = 8323;
	#10 counter$count = 8324;
	#10 counter$count = 8325;
	#10 counter$count = 8326;
	#10 counter$count = 8327;
	#10 counter$count = 8328;
	#10 counter$count = 8329;
	#10 counter$count = 8330;
	#10 counter$count = 8331;
	#10 counter$count = 8332;
	#10 counter$count = 8333;
	#10 counter$count = 8334;
	#10 counter$count = 8335;
	#10 counter$count = 8336;
	#10 counter$count = 8337;
	#10 counter$count = 8338;
	#10 counter$count = 8339;
	#10 counter$count = 8340;
	#10 counter$count = 8341;
	#10 counter$count = 8342;
	#10 counter$count = 8343;
	#10 counter$count = 8344;
	#10 counter$count = 8345;
	#10 counter$count = 8346;
	#10 counter$count = 8347;
	#10 counter$count = 8348;
	#10 counter$count = 8349;
	#10 counter$count = 8350;
	#10 counter$count = 8351;
	#10 counter$count = 8352;
	#10 counter$count = 8353;
	#10 counter$count = 8354;
	#10 counter$count = 8355;
	#10 counter$count = 8356;
	#10 counter$count = 8357;
	#10 counter$count = 8358;
	#10 counter$count = 8359;
	#10 counter$count = 8360;
	#10 counter$count = 8361;
	#10 counter$count = 8362;
	#10 counter$count = 8363;
	#10 counter$count = 8364;
	#10 counter$count = 8365;
	#10 counter$count = 8366;
	#10 counter$count = 8367;
	#10 counter$count = 8368;
	#10 counter$count = 8369;
	#10 counter$count = 8370;
	#10 counter$count = 8371;
	#10 counter$count = 8372;
	#10 counter$count = 8373;
	#10 counter$count = 8374;
	#10 counter$count = 8375;
	#10 counter$count = 8376;
	#10 counter$count = 8377;
	#10 counter$count = 8378;
	#10 counter$count = 8379;
	#10 counter$count = 8380;
	#10 counter$count = 8381;
	#10 counter$count = 8382;
	#10 counter$count = 8383;
	#10 counter$count = 8384;
	#10 counter$count = 8385;
	#10 counter$count = 8386;
	#10 counter$count = 8387;
	#10 counter$count = 8388;
	#10 counter$count = 8389;
	#10 counter$count = 8390;
	#10 counter$count = 8391;
	#10 counter$count = 8392;
	#10 counter$count = 8393;
	#10 counter$count = 8394;
	#10 counter$count = 8395;
	#10 counter$count = 8396;
	#10 counter$count = 8397;
	#10 counter$count = 8398;
	#10 counter$count = 8399;
	#10 counter$count = 8400;
	#10 counter$count = 8401;
	#10 counter$count = 8402;
	#10 counter$count = 8403;
	#10 counter$count = 8404;
	#10 counter$count = 8405;
	#10 counter$count = 8406;
	#10 counter$count = 8407;
	#10 counter$count = 8408;
	#10 counter$count = 8409;
	#10 counter$count = 8410;
	#10 counter$count = 8411;
	#10 counter$count = 8412;
	#10 counter$count = 8413;
	#10 counter$count = 8414;
	#10 counter$count = 8415;
	#10 counter$count = 8416;
	#10 counter$count = 8417;
	#10 counter$count = 8418;
	#10 counter$count = 8419;
	#10 counter$count = 8420;
	#10 counter$count = 8421;
	#10 counter$count = 8422;
	#10 counter$count = 8423;
	#10 counter$count = 8424;
	#10 counter$count = 8425;
	#10 counter$count = 8426;
	#10 counter$count = 8427;
	#10 counter$count = 8428;
	#10 counter$count = 8429;
	#10 counter$count = 8430;
	#10 counter$count = 8431;
	#10 counter$count = 8432;
	#10 counter$count = 8433;
	#10 counter$count = 8434;
	#10 counter$count = 8435;
	#10 counter$count = 8436;
	#10 counter$count = 8437;
	#10 counter$count = 8438;
	#10 counter$count = 8439;
	#10 counter$count = 8440;
	#10 counter$count = 8441;
	#10 counter$count = 8442;
	#10 counter$count = 8443;
	#10 counter$count = 8444;
	#10 counter$count = 8445;
	#10 counter$count = 8446;
	#10 counter$count = 8447;
	#10 counter$count = 8448;
	#10 counter$count = 8449;
	#10 counter$count = 8450;
	#10 counter$count = 8451;
	#10 counter$count = 8452;
	#10 counter$count = 8453;
	#10 counter$count = 8454;
	#10 counter$count = 8455;
	#10 counter$count = 8456;
	#10 counter$count = 8457;
	#10 counter$count = 8458;
	#10 counter$count = 8459;
	#10 counter$count = 8460;
	#10 counter$count = 8461;
	#10 counter$count = 8462;
	#10 counter$count = 8463;
	#10 counter$count = 8464;
	#10 counter$count = 8465;
	#10 counter$count = 8466;
	#10 counter$count = 8467;
	#10 counter$count = 8468;
	#10 counter$count = 8469;
	#10 counter$count = 8470;
	#10 counter$count = 8471;
	#10 counter$count = 8472;
	#10 counter$count = 8473;
	#10 counter$count = 8474;
	#10 counter$count = 8475;
	#10 counter$count = 8476;
	#10 counter$count = 8477;
	#10 counter$count = 8478;
	#10 counter$count = 8479;
	#10 counter$count = 8480;
	#10 counter$count = 8481;
	#10 counter$count = 8482;
	#10 counter$count = 8483;
	#10 counter$count = 8484;
	#10 counter$count = 8485;
	#10 counter$count = 8486;
	#10 counter$count = 8487;
	#10 counter$count = 8488;
	#10 counter$count = 8489;
	#10 counter$count = 8490;
	#10 counter$count = 8491;
	#10 counter$count = 8492;
	#10 counter$count = 8493;
	#10 counter$count = 8494;
	#10 counter$count = 8495;
	#10 counter$count = 8496;
	#10 counter$count = 8497;
	#10 counter$count = 8498;
	#10 counter$count = 8499;
	#10 counter$count = 8500;
	#10 counter$count = 8501;
	#10 counter$count = 8502;
	#10 counter$count = 8503;
	#10 counter$count = 8504;
	#10 counter$count = 8505;
	#10 counter$count = 8506;
	#10 counter$count = 8507;
	#10 counter$count = 8508;
	#10 counter$count = 8509;
	#10 counter$count = 8510;
	#10 counter$count = 8511;
	#10 counter$count = 8512;
	#10 counter$count = 8513;
	#10 counter$count = 8514;
	#10 counter$count = 8515;
	#10 counter$count = 8516;
	#10 counter$count = 8517;
	#10 counter$count = 8518;
	#10 counter$count = 8519;
	#10 counter$count = 8520;
	#10 counter$count = 8521;
	#10 counter$count = 8522;
	#10 counter$count = 8523;
	#10 counter$count = 8524;
	#10 counter$count = 8525;
	#10 counter$count = 8526;
	#10 counter$count = 8527;
	#10 counter$count = 8528;
	#10 counter$count = 8529;
	#10 counter$count = 8530;
	#10 counter$count = 8531;
	#10 counter$count = 8532;
	#10 counter$count = 8533;
	#10 counter$count = 8534;
	#10 counter$count = 8535;
	#10 counter$count = 8536;
	#10 counter$count = 8537;
	#10 counter$count = 8538;
	#10 counter$count = 8539;
	#10 counter$count = 8540;
	#10 counter$count = 8541;
	#10 counter$count = 8542;
	#10 counter$count = 8543;
	#10 counter$count = 8544;
	#10 counter$count = 8545;
	#10 counter$count = 8546;
	#10 counter$count = 8547;
	#10 counter$count = 8548;
	#10 counter$count = 8549;
	#10 counter$count = 8550;
	#10 counter$count = 8551;
	#10 counter$count = 8552;
	#10 counter$count = 8553;
	#10 counter$count = 8554;
	#10 counter$count = 8555;
	#10 counter$count = 8556;
	#10 counter$count = 8557;
	#10 counter$count = 8558;
	#10 counter$count = 8559;
	#10 counter$count = 8560;
	#10 counter$count = 8561;
	#10 counter$count = 8562;
	#10 counter$count = 8563;
	#10 counter$count = 8564;
	#10 counter$count = 8565;
	#10 counter$count = 8566;
	#10 counter$count = 8567;
	#10 counter$count = 8568;
	#10 counter$count = 8569;
	#10 counter$count = 8570;
	#10 counter$count = 8571;
	#10 counter$count = 8572;
	#10 counter$count = 8573;
	#10 counter$count = 8574;
	#10 counter$count = 8575;
	#10 counter$count = 8576;
	#10 counter$count = 8577;
	#10 counter$count = 8578;
	#10 counter$count = 8579;
	#10 counter$count = 8580;
	#10 counter$count = 8581;
	#10 counter$count = 8582;
	#10 counter$count = 8583;
	#10 counter$count = 8584;
	#10 counter$count = 8585;
	#10 counter$count = 8586;
	#10 counter$count = 8587;
	#10 counter$count = 8588;
	#10 counter$count = 8589;
	#10 counter$count = 8590;
	#10 counter$count = 8591;
	#10 counter$count = 8592;
	#10 counter$count = 8593;
	#10 counter$count = 8594;
	#10 counter$count = 8595;
	#10 counter$count = 8596;
	#10 counter$count = 8597;
	#10 counter$count = 8598;
	#10 counter$count = 8599;
	#10 counter$count = 8600;
	#10 counter$count = 8601;
	#10 counter$count = 8602;
	#10 counter$count = 8603;
	#10 counter$count = 8604;
	#10 counter$count = 8605;
	#10 counter$count = 8606;
	#10 counter$count = 8607;
	#10 counter$count = 8608;
	#10 counter$count = 8609;
	#10 counter$count = 8610;
	#10 counter$count = 8611;
	#10 counter$count = 8612;
	#10 counter$count = 8613;
	#10 counter$count = 8614;
	#10 counter$count = 8615;
	#10 counter$count = 8616;
	#10 counter$count = 8617;
	#10 counter$count = 8618;
	#10 counter$count = 8619;
	#10 counter$count = 8620;
	#10 counter$count = 8621;
	#10 counter$count = 8622;
	#10 counter$count = 8623;
	#10 counter$count = 8624;
	#10 counter$count = 8625;
	#10 counter$count = 8626;
	#10 counter$count = 8627;
	#10 counter$count = 8628;
	#10 counter$count = 8629;
	#10 counter$count = 8630;
	#10 counter$count = 8631;
	#10 counter$count = 8632;
	#10 counter$count = 8633;
	#10 counter$count = 8634;
	#10 counter$count = 8635;
	#10 counter$count = 8636;
	#10 counter$count = 8637;
	#10 counter$count = 8638;
	#10 counter$count = 8639;
	#10 counter$count = 8640;
	#10 counter$count = 8641;
	#10 counter$count = 8642;
	#10 counter$count = 8643;
	#10 counter$count = 8644;
	#10 counter$count = 8645;
	#10 counter$count = 8646;
	#10 counter$count = 8647;
	#10 counter$count = 8648;
	#10 counter$count = 8649;
	#10 counter$count = 8650;
	#10 counter$count = 8651;
	#10 counter$count = 8652;
	#10 counter$count = 8653;
	#10 counter$count = 8654;
	#10 counter$count = 8655;
	#10 counter$count = 8656;
	#10 counter$count = 8657;
	#10 counter$count = 8658;
	#10 counter$count = 8659;
	#10 counter$count = 8660;
	#10 counter$count = 8661;
	#10 counter$count = 8662;
	#10 counter$count = 8663;
	#10 counter$count = 8664;
	#10 counter$count = 8665;
	#10 counter$count = 8666;
	#10 counter$count = 8667;
	#10 counter$count = 8668;
	#10 counter$count = 8669;
	#10 counter$count = 8670;
	#10 counter$count = 8671;
	#10 counter$count = 8672;
	#10 counter$count = 8673;
	#10 counter$count = 8674;
	#10 counter$count = 8675;
	#10 counter$count = 8676;
	#10 counter$count = 8677;
	#10 counter$count = 8678;
	#10 counter$count = 8679;
	#10 counter$count = 8680;
	#10 counter$count = 8681;
	#10 counter$count = 8682;
	#10 counter$count = 8683;
	#10 counter$count = 8684;
	#10 counter$count = 8685;
	#10 counter$count = 8686;
	#10 counter$count = 8687;
	#10 counter$count = 8688;
	#10 counter$count = 8689;
	#10 counter$count = 8690;
	#10 counter$count = 8691;
	#10 counter$count = 8692;
	#10 counter$count = 8693;
	#10 counter$count = 8694;
	#10 counter$count = 8695;
	#10 counter$count = 8696;
	#10 counter$count = 8697;
	#10 counter$count = 8698;
	#10 counter$count = 8699;
	#10 counter$count = 8700;
	#10 counter$count = 8701;
	#10 counter$count = 8702;
	#10 counter$count = 8703;
	#10 counter$count = 8704;
	#10 counter$count = 8705;
	#10 counter$count = 8706;
	#10 counter$count = 8707;
	#10 counter$count = 8708;
	#10 counter$count = 8709;
	#10 counter$count = 8710;
	#10 counter$count = 8711;
	#10 counter$count = 8712;
	#10 counter$count = 8713;
	#10 counter$count = 8714;
	#10 counter$count = 8715;
	#10 counter$count = 8716;
	#10 counter$count = 8717;
	#10 counter$count = 8718;
	#10 counter$count = 8719;
	#10 counter$count = 8720;
	#10 counter$count = 8721;
	#10 counter$count = 8722;
	#10 counter$count = 8723;
	#10 counter$count = 8724;
	#10 counter$count = 8725;
	#10 counter$count = 8726;
	#10 counter$count = 8727;
	#10 counter$count = 8728;
	#10 counter$count = 8729;
	#10 counter$count = 8730;
	#10 counter$count = 8731;
	#10 counter$count = 8732;
	#10 counter$count = 8733;
	#10 counter$count = 8734;
	#10 counter$count = 8735;
	#10 counter$count = 8736;
	#10 counter$count = 8737;
	#10 counter$count = 8738;
	#10 counter$count = 8739;
	#10 counter$count = 8740;
	#10 counter$count = 8741;
	#10 counter$count = 8742;
	#10 counter$count = 8743;
	#10 counter$count = 8744;
	#10 counter$count = 8745;
	#10 counter$count = 8746;
	#10 counter$count = 8747;
	#10 counter$count = 8748;
	#10 counter$count = 8749;
	#10 counter$count = 8750;
	#10 counter$count = 8751;
	#10 counter$count = 8752;
	#10 counter$count = 8753;
	#10 counter$count = 8754;
	#10 counter$count = 8755;
	#10 counter$count = 8756;
	#10 counter$count = 8757;
	#10 counter$count = 8758;
	#10 counter$count = 8759;
	#10 counter$count = 8760;
	#10 counter$count = 8761;
	#10 counter$count = 8762;
	#10 counter$count = 8763;
	#10 counter$count = 8764;
	#10 counter$count = 8765;
	#10 counter$count = 8766;
	#10 counter$count = 8767;
	#10 counter$count = 8768;
	#10 counter$count = 8769;
	#10 counter$count = 8770;
	#10 counter$count = 8771;
	#10 counter$count = 8772;
	#10 counter$count = 8773;
	#10 counter$count = 8774;
	#10 counter$count = 8775;
	#10 counter$count = 8776;
	#10 counter$count = 8777;
	#10 counter$count = 8778;
	#10 counter$count = 8779;
	#10 counter$count = 8780;
	#10 counter$count = 8781;
	#10 counter$count = 8782;
	#10 counter$count = 8783;
	#10 counter$count = 8784;
	#10 counter$count = 8785;
	#10 counter$count = 8786;
	#10 counter$count = 8787;
	#10 counter$count = 8788;
	#10 counter$count = 8789;
	#10 counter$count = 8790;
	#10 counter$count = 8791;
	#10 counter$count = 8792;
	#10 counter$count = 8793;
	#10 counter$count = 8794;
	#10 counter$count = 8795;
	#10 counter$count = 8796;
	#10 counter$count = 8797;
	#10 counter$count = 8798;
	#10 counter$count = 8799;
	#10 counter$count = 8800;
	#10 counter$count = 8801;
	#10 counter$count = 8802;
	#10 counter$count = 8803;
	#10 counter$count = 8804;
	#10 counter$count = 8805;
	#10 counter$count = 8806;
	#10 counter$count = 8807;
	#10 counter$count = 8808;
	#10 counter$count = 8809;
	#10 counter$count = 8810;
	#10 counter$count = 8811;
	#10 counter$count = 8812;
	#10 counter$count = 8813;
	#10 counter$count = 8814;
	#10 counter$count = 8815;
	#10 counter$count = 8816;
	#10 counter$count = 8817;
	#10 counter$count = 8818;
	#10 counter$count = 8819;
	#10 counter$count = 8820;
	#10 counter$count = 8821;
	#10 counter$count = 8822;
	#10 counter$count = 8823;
	#10 counter$count = 8824;
	#10 counter$count = 8825;
	#10 counter$count = 8826;
	#10 counter$count = 8827;
	#10 counter$count = 8828;
	#10 counter$count = 8829;
	#10 counter$count = 8830;
	#10 counter$count = 8831;
	#10 counter$count = 8832;
	#10 counter$count = 8833;
	#10 counter$count = 8834;
	#10 counter$count = 8835;
	#10 counter$count = 8836;
	#10 counter$count = 8837;
	#10 counter$count = 8838;
	#10 counter$count = 8839;
	#10 counter$count = 8840;
	#10 counter$count = 8841;
	#10 counter$count = 8842;
	#10 counter$count = 8843;
	#10 counter$count = 8844;
	#10 counter$count = 8845;
	#10 counter$count = 8846;
	#10 counter$count = 8847;
	#10 counter$count = 8848;
	#10 counter$count = 8849;
	#10 counter$count = 8850;
	#10 counter$count = 8851;
	#10 counter$count = 8852;
	#10 counter$count = 8853;
	#10 counter$count = 8854;
	#10 counter$count = 8855;
	#10 counter$count = 8856;
	#10 counter$count = 8857;
	#10 counter$count = 8858;
	#10 counter$count = 8859;
	#10 counter$count = 8860;
	#10 counter$count = 8861;
	#10 counter$count = 8862;
	#10 counter$count = 8863;
	#10 counter$count = 8864;
	#10 counter$count = 8865;
	#10 counter$count = 8866;
	#10 counter$count = 8867;
	#10 counter$count = 8868;
	#10 counter$count = 8869;
	#10 counter$count = 8870;
	#10 counter$count = 8871;
	#10 counter$count = 8872;
	#10 counter$count = 8873;
	#10 counter$count = 8874;
	#10 counter$count = 8875;
	#10 counter$count = 8876;
	#10 counter$count = 8877;
	#10 counter$count = 8878;
	#10 counter$count = 8879;
	#10 counter$count = 8880;
	#10 counter$count = 8881;
	#10 counter$count = 8882;
	#10 counter$count = 8883;
	#10 counter$count = 8884;
	#10 counter$count = 8885;
	#10 counter$count = 8886;
	#10 counter$count = 8887;
	#10 counter$count = 8888;
	#10 counter$count = 8889;
	#10 counter$count = 8890;
	#10 counter$count = 8891;
	#10 counter$count = 8892;
	#10 counter$count = 8893;
	#10 counter$count = 8894;
	#10 counter$count = 8895;
	#10 counter$count = 8896;
	#10 counter$count = 8897;
	#10 counter$count = 8898;
	#10 counter$count = 8899;
	#10 counter$count = 8900;
	#10 counter$count = 8901;
	#10 counter$count = 8902;
	#10 counter$count = 8903;
	#10 counter$count = 8904;
	#10 counter$count = 8905;
	#10 counter$count = 8906;
	#10 counter$count = 8907;
	#10 counter$count = 8908;
	#10 counter$count = 8909;
	#10 counter$count = 8910;
	#10 counter$count = 8911;
	#10 counter$count = 8912;
	#10 counter$count = 8913;
	#10 counter$count = 8914;
	#10 counter$count = 8915;
	#10 counter$count = 8916;
	#10 counter$count = 8917;
	#10 counter$count = 8918;
	#10 counter$count = 8919;
	#10 counter$count = 8920;
	#10 counter$count = 8921;
	#10 counter$count = 8922;
	#10 counter$count = 8923;
	#10 counter$count = 8924;
	#10 counter$count = 8925;
	#10 counter$count = 8926;
	#10 counter$count = 8927;
	#10 counter$count = 8928;
	#10 counter$count = 8929;
	#10 counter$count = 8930;
	#10 counter$count = 8931;
	#10 counter$count = 8932;
	#10 counter$count = 8933;
	#10 counter$count = 8934;
	#10 counter$count = 8935;
	#10 counter$count = 8936;
	#10 counter$count = 8937;
	#10 counter$count = 8938;
	#10 counter$count = 8939;
	#10 counter$count = 8940;
	#10 counter$count = 8941;
	#10 counter$count = 8942;
	#10 counter$count = 8943;
	#10 counter$count = 8944;
	#10 counter$count = 8945;
	#10 counter$count = 8946;
	#10 counter$count = 8947;
	#10 counter$count = 8948;
	#10 counter$count = 8949;
	#10 counter$count = 8950;
	#10 counter$count = 8951;
	#10 counter$count = 8952;
	#10 counter$count = 8953;
	#10 counter$count = 8954;
	#10 counter$count = 8955;
	#10 counter$count = 8956;
	#10 counter$count = 8957;
	#10 counter$count = 8958;
	#10 counter$count = 8959;
	#10 counter$count = 8960;
	#10 counter$count = 8961;
	#10 counter$count = 8962;
	#10 counter$count = 8963;
	#10 counter$count = 8964;
	#10 counter$count = 8965;
	#10 counter$count = 8966;
	#10 counter$count = 8967;
	#10 counter$count = 8968;
	#10 counter$count = 8969;
	#10 counter$count = 8970;
	#10 counter$count = 8971;
	#10 counter$count = 8972;
	#10 counter$count = 8973;
	#10 counter$count = 8974;
	#10 counter$count = 8975;
	#10 counter$count = 8976;
	#10 counter$count = 8977;
	#10 counter$count = 8978;
	#10 counter$count = 8979;
	#10 counter$count = 8980;
	#10 counter$count = 8981;
	#10 counter$count = 8982;
	#10 counter$count = 8983;
	#10 counter$count = 8984;
	#10 counter$count = 8985;
	#10 counter$count = 8986;
	#10 counter$count = 8987;
	#10 counter$count = 8988;
	#10 counter$count = 8989;
	#10 counter$count = 8990;
	#10 counter$count = 8991;
	#10 counter$count = 8992;
	#10 counter$count = 8993;
	#10 counter$count = 8994;
	#10 counter$count = 8995;
	#10 counter$count = 8996;
	#10 counter$count = 8997;
	#10 counter$count = 8998;
	#10 counter$count = 8999;
	#10 counter$count = 9000;
	#10 counter$count = 9001;
	#10 counter$count = 9002;
	#10 counter$count = 9003;
	#10 counter$count = 9004;
	#10 counter$count = 9005;
	#10 counter$count = 9006;
	#10 counter$count = 9007;
	#10 counter$count = 9008;
	#10 counter$count = 9009;
	#10 counter$count = 9010;
	#10 counter$count = 9011;
	#10 counter$count = 9012;
	#10 counter$count = 9013;
	#10 counter$count = 9014;
	#10 counter$count = 9015;
	#10 counter$count = 9016;
	#10 counter$count = 9017;
	#10 counter$count = 9018;
	#10 counter$count = 9019;
	#10 counter$count = 9020;
	#10 counter$count = 9021;
	#10 counter$count = 9022;
	#10 counter$count = 9023;
	#10 counter$count = 9024;
	#10 counter$count = 9025;
	#10 counter$count = 9026;
	#10 counter$count = 9027;
	#10 counter$count = 9028;
	#10 counter$count = 9029;
	#10 counter$count = 9030;
	#10 counter$count = 9031;
	#10 counter$count = 9032;
	#10 counter$count = 9033;
	#10 counter$count = 9034;
	#10 counter$count = 9035;
	#10 counter$count = 9036;
	#10 counter$count = 9037;
	#10 counter$count = 9038;
	#10 counter$count = 9039;
	#10 counter$count = 9040;
	#10 counter$count = 9041;
	#10 counter$count = 9042;
	#10 counter$count = 9043;
	#10 counter$count = 9044;
	#10 counter$count = 9045;
	#10 counter$count = 9046;
	#10 counter$count = 9047;
	#10 counter$count = 9048;
	#10 counter$count = 9049;
	#10 counter$count = 9050;
	#10 counter$count = 9051;
	#10 counter$count = 9052;
	#10 counter$count = 9053;
	#10 counter$count = 9054;
	#10 counter$count = 9055;
	#10 counter$count = 9056;
	#10 counter$count = 9057;
	#10 counter$count = 9058;
	#10 counter$count = 9059;
	#10 counter$count = 9060;
	#10 counter$count = 9061;
	#10 counter$count = 9062;
	#10 counter$count = 9063;
	#10 counter$count = 9064;
	#10 counter$count = 9065;
	#10 counter$count = 9066;
	#10 counter$count = 9067;
	#10 counter$count = 9068;
	#10 counter$count = 9069;
	#10 counter$count = 9070;
	#10 counter$count = 9071;
	#10 counter$count = 9072;
	#10 counter$count = 9073;
	#10 counter$count = 9074;
	#10 counter$count = 9075;
	#10 counter$count = 9076;
	#10 counter$count = 9077;
	#10 counter$count = 9078;
	#10 counter$count = 9079;
	#10 counter$count = 9080;
	#10 counter$count = 9081;
	#10 counter$count = 9082;
	#10 counter$count = 9083;
	#10 counter$count = 9084;
	#10 counter$count = 9085;
	#10 counter$count = 9086;
	#10 counter$count = 9087;
	#10 counter$count = 9088;
	#10 counter$count = 9089;
	#10 counter$count = 9090;
	#10 counter$count = 9091;
	#10 counter$count = 9092;
	#10 counter$count = 9093;
	#10 counter$count = 9094;
	#10 counter$count = 9095;
	#10 counter$count = 9096;
	#10 counter$count = 9097;
	#10 counter$count = 9098;
	#10 counter$count = 9099;
	#10 counter$count = 9100;
	#10 counter$count = 9101;
	#10 counter$count = 9102;
	#10 counter$count = 9103;
	#10 counter$count = 9104;
	#10 counter$count = 9105;
	#10 counter$count = 9106;
	#10 counter$count = 9107;
	#10 counter$count = 9108;
	#10 counter$count = 9109;
	#10 counter$count = 9110;
	#10 counter$count = 9111;
	#10 counter$count = 9112;
	#10 counter$count = 9113;
	#10 counter$count = 9114;
	#10 counter$count = 9115;
	#10 counter$count = 9116;
	#10 counter$count = 9117;
	#10 counter$count = 9118;
	#10 counter$count = 9119;
	#10 counter$count = 9120;
	#10 counter$count = 9121;
	#10 counter$count = 9122;
	#10 counter$count = 9123;
	#10 counter$count = 9124;
	#10 counter$count = 9125;
	#10 counter$count = 9126;
	#10 counter$count = 9127;
	#10 counter$count = 9128;
	#10 counter$count = 9129;
	#10 counter$count = 9130;
	#10 counter$count = 9131;
	#10 counter$count = 9132;
	#10 counter$count = 9133;
	#10 counter$count = 9134;
	#10 counter$count = 9135;
	#10 counter$count = 9136;
	#10 counter$count = 9137;
	#10 counter$count = 9138;
	#10 counter$count = 9139;
	#10 counter$count = 9140;
	#10 counter$count = 9141;
	#10 counter$count = 9142;
	#10 counter$count = 9143;
	#10 counter$count = 9144;
	#10 counter$count = 9145;
	#10 counter$count = 9146;
	#10 counter$count = 9147;
	#10 counter$count = 9148;
	#10 counter$count = 9149;
	#10 counter$count = 9150;
	#10 counter$count = 9151;
	#10 counter$count = 9152;
	#10 counter$count = 9153;
	#10 counter$count = 9154;
	#10 counter$count = 9155;
	#10 counter$count = 9156;
	#10 counter$count = 9157;
	#10 counter$count = 9158;
	#10 counter$count = 9159;
	#10 counter$count = 9160;
	#10 counter$count = 9161;
	#10 counter$count = 9162;
	#10 counter$count = 9163;
	#10 counter$count = 9164;
	#10 counter$count = 9165;
	#10 counter$count = 9166;
	#10 counter$count = 9167;
	#10 counter$count = 9168;
	#10 counter$count = 9169;
	#10 counter$count = 9170;
	#10 counter$count = 9171;
	#10 counter$count = 9172;
	#10 counter$count = 9173;
	#10 counter$count = 9174;
	#10 counter$count = 9175;
	#10 counter$count = 9176;
	#10 counter$count = 9177;
	#10 counter$count = 9178;
	#10 counter$count = 9179;
	#10 counter$count = 9180;
	#10 counter$count = 9181;
	#10 counter$count = 9182;
	#10 counter$count = 9183;
	#10 counter$count = 9184;
	#10 counter$count = 9185;
	#10 counter$count = 9186;
	#10 counter$count = 9187;
	#10 counter$count = 9188;
	#10 counter$count = 9189;
	#10 counter$count = 9190;
	#10 counter$count = 9191;
	#10 counter$count = 9192;
	#10 counter$count = 9193;
	#10 counter$count = 9194;
	#10 counter$count = 9195;
	#10 counter$count = 9196;
	#10 counter$count = 9197;
	#10 counter$count = 9198;
	#10 counter$count = 9199;
	#10 counter$count = 9200;
	#10 counter$count = 9201;
	#10 counter$count = 9202;
	#10 counter$count = 9203;
	#10 counter$count = 9204;
	#10 counter$count = 9205;
	#10 counter$count = 9206;
	#10 counter$count = 9207;
	#10 counter$count = 9208;
	#10 counter$count = 9209;
	#10 counter$count = 9210;
	#10 counter$count = 9211;
	#10 counter$count = 9212;
	#10 counter$count = 9213;
	#10 counter$count = 9214;
	#10 counter$count = 9215;
	#10 counter$count = 9216;
	#10 counter$count = 9217;
	#10 counter$count = 9218;
	#10 counter$count = 9219;
	#10 counter$count = 9220;
	#10 counter$count = 9221;
	#10 counter$count = 9222;
	#10 counter$count = 9223;
	#10 counter$count = 9224;
	#10 counter$count = 9225;
	#10 counter$count = 9226;
	#10 counter$count = 9227;
	#10 counter$count = 9228;
	#10 counter$count = 9229;
	#10 counter$count = 9230;
	#10 counter$count = 9231;
	#10 counter$count = 9232;
	#10 counter$count = 9233;
	#10 counter$count = 9234;
	#10 counter$count = 9235;
	#10 counter$count = 9236;
	#10 counter$count = 9237;
	#10 counter$count = 9238;
	#10 counter$count = 9239;
	#10 counter$count = 9240;
	#10 counter$count = 9241;
	#10 counter$count = 9242;
	#10 counter$count = 9243;
	#10 counter$count = 9244;
	#10 counter$count = 9245;
	#10 counter$count = 9246;
	#10 counter$count = 9247;
	#10 counter$count = 9248;
	#10 counter$count = 9249;
	#10 counter$count = 9250;
	#10 counter$count = 9251;
	#10 counter$count = 9252;
	#10 counter$count = 9253;
	#10 counter$count = 9254;
	#10 counter$count = 9255;
	#10 counter$count = 9256;
	#10 counter$count = 9257;
	#10 counter$count = 9258;
	#10 counter$count = 9259;
	#10 counter$count = 9260;
	#10 counter$count = 9261;
	#10 counter$count = 9262;
	#10 counter$count = 9263;
	#10 counter$count = 9264;
	#10 counter$count = 9265;
	#10 counter$count = 9266;
	#10 counter$count = 9267;
	#10 counter$count = 9268;
	#10 counter$count = 9269;
	#10 counter$count = 9270;
	#10 counter$count = 9271;
	#10 counter$count = 9272;
	#10 counter$count = 9273;
	#10 counter$count = 9274;
	#10 counter$count = 9275;
	#10 counter$count = 9276;
	#10 counter$count = 9277;
	#10 counter$count = 9278;
	#10 counter$count = 9279;
	#10 counter$count = 9280;
	#10 counter$count = 9281;
	#10 counter$count = 9282;
	#10 counter$count = 9283;
	#10 counter$count = 9284;
	#10 counter$count = 9285;
	#10 counter$count = 9286;
	#10 counter$count = 9287;
	#10 counter$count = 9288;
	#10 counter$count = 9289;
	#10 counter$count = 9290;
	#10 counter$count = 9291;
	#10 counter$count = 9292;
	#10 counter$count = 9293;
	#10 counter$count = 9294;
	#10 counter$count = 9295;
	#10 counter$count = 9296;
	#10 counter$count = 9297;
	#10 counter$count = 9298;
	#10 counter$count = 9299;
	#10 counter$count = 9300;
	#10 counter$count = 9301;
	#10 counter$count = 9302;
	#10 counter$count = 9303;
	#10 counter$count = 9304;
	#10 counter$count = 9305;
	#10 counter$count = 9306;
	#10 counter$count = 9307;
	#10 counter$count = 9308;
	#10 counter$count = 9309;
	#10 counter$count = 9310;
	#10 counter$count = 9311;
	#10 counter$count = 9312;
	#10 counter$count = 9313;
	#10 counter$count = 9314;
	#10 counter$count = 9315;
	#10 counter$count = 9316;
	#10 counter$count = 9317;
	#10 counter$count = 9318;
	#10 counter$count = 9319;
	#10 counter$count = 9320;
	#10 counter$count = 9321;
	#10 counter$count = 9322;
	#10 counter$count = 9323;
	#10 counter$count = 9324;
	#10 counter$count = 9325;
	#10 counter$count = 9326;
	#10 counter$count = 9327;
	#10 counter$count = 9328;
	#10 counter$count = 9329;
	#10 counter$count = 9330;
	#10 counter$count = 9331;
	#10 counter$count = 9332;
	#10 counter$count = 9333;
	#10 counter$count = 9334;
	#10 counter$count = 9335;
	#10 counter$count = 9336;
	#10 counter$count = 9337;
	#10 counter$count = 9338;
	#10 counter$count = 9339;
	#10 counter$count = 9340;
	#10 counter$count = 9341;
	#10 counter$count = 9342;
	#10 counter$count = 9343;
	#10 counter$count = 9344;
	#10 counter$count = 9345;
	#10 counter$count = 9346;
	#10 counter$count = 9347;
	#10 counter$count = 9348;
	#10 counter$count = 9349;
	#10 counter$count = 9350;
	#10 counter$count = 9351;
	#10 counter$count = 9352;
	#10 counter$count = 9353;
	#10 counter$count = 9354;
	#10 counter$count = 9355;
	#10 counter$count = 9356;
	#10 counter$count = 9357;
	#10 counter$count = 9358;
	#10 counter$count = 9359;
	#10 counter$count = 9360;
	#10 counter$count = 9361;
	#10 counter$count = 9362;
	#10 counter$count = 9363;
	#10 counter$count = 9364;
	#10 counter$count = 9365;
	#10 counter$count = 9366;
	#10 counter$count = 9367;
	#10 counter$count = 9368;
	#10 counter$count = 9369;
	#10 counter$count = 9370;
	#10 counter$count = 9371;
	#10 counter$count = 9372;
	#10 counter$count = 9373;
	#10 counter$count = 9374;
	#10 counter$count = 9375;
	#10 counter$count = 9376;
	#10 counter$count = 9377;
	#10 counter$count = 9378;
	#10 counter$count = 9379;
	#10 counter$count = 9380;
	#10 counter$count = 9381;
	#10 counter$count = 9382;
	#10 counter$count = 9383;
	#10 counter$count = 9384;
	#10 counter$count = 9385;
	#10 counter$count = 9386;
	#10 counter$count = 9387;
	#10 counter$count = 9388;
	#10 counter$count = 9389;
	#10 counter$count = 9390;
	#10 counter$count = 9391;
	#10 counter$count = 9392;
	#10 counter$count = 9393;
	#10 counter$count = 9394;
	#10 counter$count = 9395;
	#10 counter$count = 9396;
	#10 counter$count = 9397;
	#10 counter$count = 9398;
	#10 counter$count = 9399;
	#10 counter$count = 9400;
	#10 counter$count = 9401;
	#10 counter$count = 9402;
	#10 counter$count = 9403;
	#10 counter$count = 9404;
	#10 counter$count = 9405;
	#10 counter$count = 9406;
	#10 counter$count = 9407;
	#10 counter$count = 9408;
	#10 counter$count = 9409;
	#10 counter$count = 9410;
	#10 counter$count = 9411;
	#10 counter$count = 9412;
	#10 counter$count = 9413;
	#10 counter$count = 9414;
	#10 counter$count = 9415;
	#10 counter$count = 9416;
	#10 counter$count = 9417;
	#10 counter$count = 9418;
	#10 counter$count = 9419;
	#10 counter$count = 9420;
	#10 counter$count = 9421;
	#10 counter$count = 9422;
	#10 counter$count = 9423;
	#10 counter$count = 9424;
	#10 counter$count = 9425;
	#10 counter$count = 9426;
	#10 counter$count = 9427;
	#10 counter$count = 9428;
	#10 counter$count = 9429;
	#10 counter$count = 9430;
	#10 counter$count = 9431;
	#10 counter$count = 9432;
	#10 counter$count = 9433;
	#10 counter$count = 9434;
	#10 counter$count = 9435;
	#10 counter$count = 9436;
	#10 counter$count = 9437;
	#10 counter$count = 9438;
	#10 counter$count = 9439;
	#10 counter$count = 9440;
	#10 counter$count = 9441;
	#10 counter$count = 9442;
	#10 counter$count = 9443;
	#10 counter$count = 9444;
	#10 counter$count = 9445;
	#10 counter$count = 9446;
	#10 counter$count = 9447;
	#10 counter$count = 9448;
	#10 counter$count = 9449;
	#10 counter$count = 9450;
	#10 counter$count = 9451;
	#10 counter$count = 9452;
	#10 counter$count = 9453;
	#10 counter$count = 9454;
	#10 counter$count = 9455;
	#10 counter$count = 9456;
	#10 counter$count = 9457;
	#10 counter$count = 9458;
	#10 counter$count = 9459;
	#10 counter$count = 9460;
	#10 counter$count = 9461;
	#10 counter$count = 9462;
	#10 counter$count = 9463;
	#10 counter$count = 9464;
	#10 counter$count = 9465;
	#10 counter$count = 9466;
	#10 counter$count = 9467;
	#10 counter$count = 9468;
	#10 counter$count = 9469;
	#10 counter$count = 9470;
	#10 counter$count = 9471;
	#10 counter$count = 9472;
	#10 counter$count = 9473;
	#10 counter$count = 9474;
	#10 counter$count = 9475;
	#10 counter$count = 9476;
	#10 counter$count = 9477;
	#10 counter$count = 9478;
	#10 counter$count = 9479;
	#10 counter$count = 9480;
	#10 counter$count = 9481;
	#10 counter$count = 9482;
	#10 counter$count = 9483;
	#10 counter$count = 9484;
	#10 counter$count = 9485;
	#10 counter$count = 9486;
	#10 counter$count = 9487;
	#10 counter$count = 9488;
	#10 counter$count = 9489;
	#10 counter$count = 9490;
	#10 counter$count = 9491;
	#10 counter$count = 9492;
	#10 counter$count = 9493;
	#10 counter$count = 9494;
	#10 counter$count = 9495;
	#10 counter$count = 9496;
	#10 counter$count = 9497;
	#10 counter$count = 9498;
	#10 counter$count = 9499;
	#10 counter$count = 9500;
	#10 counter$count = 9501;
	#10 counter$count = 9502;
	#10 counter$count = 9503;
	#10 counter$count = 9504;
	#10 counter$count = 9505;
	#10 counter$count = 9506;
	#10 counter$count = 9507;
	#10 counter$count = 9508;
	#10 counter$count = 9509;
	#10 counter$count = 9510;
	#10 counter$count = 9511;
	#10 counter$count = 9512;
	#10 counter$count = 9513;
	#10 counter$count = 9514;
	#10 counter$count = 9515;
	#10 counter$count = 9516;
	#10 counter$count = 9517;
	#10 counter$count = 9518;
	#10 counter$count = 9519;
	#10 counter$count = 9520;
	#10 counter$count = 9521;
	#10 counter$count = 9522;
	#10 counter$count = 9523;
	#10 counter$count = 9524;
	#10 counter$count = 9525;
	#10 counter$count = 9526;
	#10 counter$count = 9527;
	#10 counter$count = 9528;
	#10 counter$count = 9529;
	#10 counter$count = 9530;
	#10 counter$count = 9531;
	#10 counter$count = 9532;
	#10 counter$count = 9533;
	#10 counter$count = 9534;
	#10 counter$count = 9535;
	#10 counter$count = 9536;
	#10 counter$count = 9537;
	#10 counter$count = 9538;
	#10 counter$count = 9539;
	#10 counter$count = 9540;
	#10 counter$count = 9541;
	#10 counter$count = 9542;
	#10 counter$count = 9543;
	#10 counter$count = 9544;
	#10 counter$count = 9545;
	#10 counter$count = 9546;
	#10 counter$count = 9547;
	#10 counter$count = 9548;
	#10 counter$count = 9549;
	#10 counter$count = 9550;
	#10 counter$count = 9551;
	#10 counter$count = 9552;
	#10 counter$count = 9553;
	#10 counter$count = 9554;
	#10 counter$count = 9555;
	#10 counter$count = 9556;
	#10 counter$count = 9557;
	#10 counter$count = 9558;
	#10 counter$count = 9559;
	#10 counter$count = 9560;
	#10 counter$count = 9561;
	#10 counter$count = 9562;
	#10 counter$count = 9563;
	#10 counter$count = 9564;
	#10 counter$count = 9565;
	#10 counter$count = 9566;
	#10 counter$count = 9567;
	#10 counter$count = 9568;
	#10 counter$count = 9569;
	#10 counter$count = 9570;
	#10 counter$count = 9571;
	#10 counter$count = 9572;
	#10 counter$count = 9573;
	#10 counter$count = 9574;
	#10 counter$count = 9575;
	#10 counter$count = 9576;
	#10 counter$count = 9577;
	#10 counter$count = 9578;
	#10 counter$count = 9579;
	#10 counter$count = 9580;
	#10 counter$count = 9581;
	#10 counter$count = 9582;
	#10 counter$count = 9583;
	#10 counter$count = 9584;
	#10 counter$count = 9585;
	#10 counter$count = 9586;
	#10 counter$count = 9587;
	#10 counter$count = 9588;
	#10 counter$count = 9589;
	#10 counter$count = 9590;
	#10 counter$count = 9591;
	#10 counter$count = 9592;
	#10 counter$count = 9593;
	#10 counter$count = 9594;
	#10 counter$count = 9595;
	#10 counter$count = 9596;
	#10 counter$count = 9597;
	#10 counter$count = 9598;
	#10 counter$count = 9599;
	#10 counter$count = 9600;
	#10 counter$count = 9601;
	#10 counter$count = 9602;
	#10 counter$count = 9603;
	#10 counter$count = 9604;
	#10 counter$count = 9605;
	#10 counter$count = 9606;
	#10 counter$count = 9607;
	#10 counter$count = 9608;
	#10 counter$count = 9609;
	#10 counter$count = 9610;
	#10 counter$count = 9611;
	#10 counter$count = 9612;
	#10 counter$count = 9613;
	#10 counter$count = 9614;
	#10 counter$count = 9615;
	#10 counter$count = 9616;
	#10 counter$count = 9617;
	#10 counter$count = 9618;
	#10 counter$count = 9619;
	#10 counter$count = 9620;
	#10 counter$count = 9621;
	#10 counter$count = 9622;
	#10 counter$count = 9623;
	#10 counter$count = 9624;
	#10 counter$count = 9625;
	#10 counter$count = 9626;
	#10 counter$count = 9627;
	#10 counter$count = 9628;
	#10 counter$count = 9629;
	#10 counter$count = 9630;
	#10 counter$count = 9631;
	#10 counter$count = 9632;
	#10 counter$count = 9633;
	#10 counter$count = 9634;
	#10 counter$count = 9635;
	#10 counter$count = 9636;
	#10 counter$count = 9637;
	#10 counter$count = 9638;
	#10 counter$count = 9639;
	#10 counter$count = 9640;
	#10 counter$count = 9641;
	#10 counter$count = 9642;
	#10 counter$count = 9643;
	#10 counter$count = 9644;
	#10 counter$count = 9645;
	#10 counter$count = 9646;
	#10 counter$count = 9647;
	#10 counter$count = 9648;
	#10 counter$count = 9649;
	#10 counter$count = 9650;
	#10 counter$count = 9651;
	#10 counter$count = 9652;
	#10 counter$count = 9653;
	#10 counter$count = 9654;
	#10 counter$count = 9655;
	#10 counter$count = 9656;
	#10 counter$count = 9657;
	#10 counter$count = 9658;
	#10 counter$count = 9659;
	#10 counter$count = 9660;
	#10 counter$count = 9661;
	#10 counter$count = 9662;
	#10 counter$count = 9663;
	#10 counter$count = 9664;
	#10 counter$count = 9665;
	#10 counter$count = 9666;
	#10 counter$count = 9667;
	#10 counter$count = 9668;
	#10 counter$count = 9669;
	#10 counter$count = 9670;
	#10 counter$count = 9671;
	#10 counter$count = 9672;
	#10 counter$count = 9673;
	#10 counter$count = 9674;
	#10 counter$count = 9675;
	#10 counter$count = 9676;
	#10 counter$count = 9677;
	#10 counter$count = 9678;
	#10 counter$count = 9679;
	#10 counter$count = 9680;
	#10 counter$count = 9681;
	#10 counter$count = 9682;
	#10 counter$count = 9683;
	#10 counter$count = 9684;
	#10 counter$count = 9685;
	#10 counter$count = 9686;
	#10 counter$count = 9687;
	#10 counter$count = 9688;
	#10 counter$count = 9689;
	#10 counter$count = 9690;
	#10 counter$count = 9691;
	#10 counter$count = 9692;
	#10 counter$count = 9693;
	#10 counter$count = 9694;
	#10 counter$count = 9695;
	#10 counter$count = 9696;
	#10 counter$count = 9697;
	#10 counter$count = 9698;
	#10 counter$count = 9699;
	#10 counter$count = 9700;
	#10 counter$count = 9701;
	#10 counter$count = 9702;
	#10 counter$count = 9703;
	#10 counter$count = 9704;
	#10 counter$count = 9705;
	#10 counter$count = 9706;
	#10 counter$count = 9707;
	#10 counter$count = 9708;
	#10 counter$count = 9709;
	#10 counter$count = 9710;
	#10 counter$count = 9711;
	#10 counter$count = 9712;
	#10 counter$count = 9713;
	#10 counter$count = 9714;
	#10 counter$count = 9715;
	#10 counter$count = 9716;
	#10 counter$count = 9717;
	#10 counter$count = 9718;
	#10 counter$count = 9719;
	#10 counter$count = 9720;
	#10 counter$count = 9721;
	#10 counter$count = 9722;
	#10 counter$count = 9723;
	#10 counter$count = 9724;
	#10 counter$count = 9725;
	#10 counter$count = 9726;
	#10 counter$count = 9727;
	#10 counter$count = 9728;
	#10 counter$count = 9729;
	#10 counter$count = 9730;
	#10 counter$count = 9731;
	#10 counter$count = 9732;
	#10 counter$count = 9733;
	#10 counter$count = 9734;
	#10 counter$count = 9735;
	#10 counter$count = 9736;
	#10 counter$count = 9737;
	#10 counter$count = 9738;
	#10 counter$count = 9739;
	#10 counter$count = 9740;
	#10 counter$count = 9741;
	#10 counter$count = 9742;
	#10 counter$count = 9743;
	#10 counter$count = 9744;
	#10 counter$count = 9745;
	#10 counter$count = 9746;
	#10 counter$count = 9747;
	#10 counter$count = 9748;
	#10 counter$count = 9749;
	#10 counter$count = 9750;
	#10 counter$count = 9751;
	#10 counter$count = 9752;
	#10 counter$count = 9753;
	#10 counter$count = 9754;
	#10 counter$count = 9755;
	#10 counter$count = 9756;
	#10 counter$count = 9757;
	#10 counter$count = 9758;
	#10 counter$count = 9759;
	#10 counter$count = 9760;
	#10 counter$count = 9761;
	#10 counter$count = 9762;
	#10 counter$count = 9763;
	#10 counter$count = 9764;
	#10 counter$count = 9765;
	#10 counter$count = 9766;
	#10 counter$count = 9767;
	#10 counter$count = 9768;
	#10 counter$count = 9769;
	#10 counter$count = 9770;
	#10 counter$count = 9771;
	#10 counter$count = 9772;
	#10 counter$count = 9773;
	#10 counter$count = 9774;
	#10 counter$count = 9775;
	#10 counter$count = 9776;
	#10 counter$count = 9777;
	#10 counter$count = 9778;
	#10 counter$count = 9779;
	#10 counter$count = 9780;
	#10 counter$count = 9781;
	#10 counter$count = 9782;
	#10 counter$count = 9783;
	#10 counter$count = 9784;
	#10 counter$count = 9785;
	#10 counter$count = 9786;
	#10 counter$count = 9787;
	#10 counter$count = 9788;
	#10 counter$count = 9789;
	#10 counter$count = 9790;
	#10 counter$count = 9791;
	#10 counter$count = 9792;
	#10 counter$count = 9793;
	#10 counter$count = 9794;
	#10 counter$count = 9795;
	#10 counter$count = 9796;
	#10 counter$count = 9797;
	#10 counter$count = 9798;
	#10 counter$count = 9799;
	#10 counter$count = 9800;
	#10 counter$count = 9801;
	#10 counter$count = 9802;
	#10 counter$count = 9803;
	#10 counter$count = 9804;
	#10 counter$count = 9805;
	#10 counter$count = 9806;
	#10 counter$count = 9807;
	#10 counter$count = 9808;
	#10 counter$count = 9809;
	#10 counter$count = 9810;
	#10 counter$count = 9811;
	#10 counter$count = 9812;
	#10 counter$count = 9813;
	#10 counter$count = 9814;
	#10 counter$count = 9815;
	#10 counter$count = 9816;
	#10 counter$count = 9817;
	#10 counter$count = 9818;
	#10 counter$count = 9819;
	#10 counter$count = 9820;
	#10 counter$count = 9821;
	#10 counter$count = 9822;
	#10 counter$count = 9823;
	#10 counter$count = 9824;
	#10 counter$count = 9825;
	#10 counter$count = 9826;
	#10 counter$count = 9827;
	#10 counter$count = 9828;
	#10 counter$count = 9829;
	#10 counter$count = 9830;
	#10 counter$count = 9831;
	#10 counter$count = 9832;
	#10 counter$count = 9833;
	#10 counter$count = 9834;
	#10 counter$count = 9835;
	#10 counter$count = 9836;
	#10 counter$count = 9837;
	#10 counter$count = 9838;
	#10 counter$count = 9839;
	#10 counter$count = 9840;
	#10 counter$count = 9841;
	#10 counter$count = 9842;
	#10 counter$count = 9843;
	#10 counter$count = 9844;
	#10 counter$count = 9845;
	#10 counter$count = 9846;
	#10 counter$count = 9847;
	#10 counter$count = 9848;
	#10 counter$count = 9849;
	#10 counter$count = 9850;
	#10 counter$count = 9851;
	#10 counter$count = 9852;
	#10 counter$count = 9853;
	#10 counter$count = 9854;
	#10 counter$count = 9855;
	#10 counter$count = 9856;
	#10 counter$count = 9857;
	#10 counter$count = 9858;
	#10 counter$count = 9859;
	#10 counter$count = 9860;
	#10 counter$count = 9861;
	#10 counter$count = 9862;
	#10 counter$count = 9863;
	#10 counter$count = 9864;
	#10 counter$count = 9865;
	#10 counter$count = 9866;
	#10 counter$count = 9867;
	#10 counter$count = 9868;
	#10 counter$count = 9869;
	#10 counter$count = 9870;
	#10 counter$count = 9871;
	#10 counter$count = 9872;
	#10 counter$count = 9873;
	#10 counter$count = 9874;
	#10 counter$count = 9875;
	#10 counter$count = 9876;
	#10 counter$count = 9877;
	#10 counter$count = 9878;
	#10 counter$count = 9879;
	#10 counter$count = 9880;
	#10 counter$count = 9881;
	#10 counter$count = 9882;
	#10 counter$count = 9883;
	#10 counter$count = 9884;
	#10 counter$count = 9885;
	#10 counter$count = 9886;
	#10 counter$count = 9887;
	#10 counter$count = 9888;
	#10 counter$count = 9889;
	#10 counter$count = 9890;
	#10 counter$count = 9891;
	#10 counter$count = 9892;
	#10 counter$count = 9893;
	#10 counter$count = 9894;
	#10 counter$count = 9895;
	#10 counter$count = 9896;
	#10 counter$count = 9897;
	#10 counter$count = 9898;
	#10 counter$count = 9899;
	#10 counter$count = 9900;
	#10 counter$count = 9901;
	#10 counter$count = 9902;
	#10 counter$count = 9903;
	#10 counter$count = 9904;
	#10 counter$count = 9905;
	#10 counter$count = 9906;
	#10 counter$count = 9907;
	#10 counter$count = 9908;
	#10 counter$count = 9909;
	#10 counter$count = 9910;
	#10 counter$count = 9911;
	#10 counter$count = 9912;
	#10 counter$count = 9913;
	#10 counter$count = 9914;
	#10 counter$count = 9915;
	#10 counter$count = 9916;
	#10 counter$count = 9917;
	#10 counter$count = 9918;
	#10 counter$count = 9919;
	#10 counter$count = 9920;
	#10 counter$count = 9921;
	#10 counter$count = 9922;
	#10 counter$count = 9923;
	#10 counter$count = 9924;
	#10 counter$count = 9925;
	#10 counter$count = 9926;
	#10 counter$count = 9927;
	#10 counter$count = 9928;
	#10 counter$count = 9929;
	#10 counter$count = 9930;
	#10 counter$count = 9931;
	#10 counter$count = 9932;
	#10 counter$count = 9933;
	#10 counter$count = 9934;
	#10 counter$count = 9935;
	#10 counter$count = 9936;
	#10 counter$count = 9937;
	#10 counter$count = 9938;
	#10 counter$count = 9939;
	#10 counter$count = 9940;
	#10 counter$count = 9941;
	#10 counter$count = 9942;
	#10 counter$count = 9943;
	#10 counter$count = 9944;
	#10 counter$count = 9945;
	#10 counter$count = 9946;
	#10 counter$count = 9947;
	#10 counter$count = 9948;
	#10 counter$count = 9949;
	#10 counter$count = 9950;
	#10 counter$count = 9951;
	#10 counter$count = 9952;
	#10 counter$count = 9953;
	#10 counter$count = 9954;
	#10 counter$count = 9955;
	#10 counter$count = 9956;
	#10 counter$count = 9957;
	#10 counter$count = 9958;
	#10 counter$count = 9959;
	#10 counter$count = 9960;
	#10 counter$count = 9961;
	#10 counter$count = 9962;
	#10 counter$count = 9963;
	#10 counter$count = 9964;
	#10 counter$count = 9965;
	#10 counter$count = 9966;
	#10 counter$count = 9967;
	#10 counter$count = 9968;
	#10 counter$count = 9969;
	#10 counter$count = 9970;
	#10 counter$count = 9971;
	#10 counter$count = 9972;
	#10 counter$count = 9973;
	#10 counter$count = 9974;
	#10 counter$count = 9975;
	#10 counter$count = 9976;
	#10 counter$count = 9977;
	#10 counter$count = 9978;
	#10 counter$count = 9979;
	#10 counter$count = 9980;
	#10 counter$count = 9981;
	#10 counter$count = 9982;
	#10 counter$count = 9983;
	#10 counter$count = 9984;
	#10 counter$count = 9985;
	#10 counter$count = 9986;
	#10 counter$count = 9987;
	#10 counter$count = 9988;
	#10 counter$count = 9989;
	#10 counter$count = 9990;
	#10 counter$count = 9991;
	#10 counter$count = 9992;
	#10 counter$count = 9993;
	#10 counter$count = 9994;
	#10 counter$count = 9995;
	#10 counter$count = 9996;
	#10 counter$count = 9997;
	#10 counter$count = 9998;
	#10 counter$count = 9999;
	#10 counter$count = 10000;
	#10 counter$count = 10001;
	#10 counter$count = 10002;
	#10 counter$count = 10003;
	#10 counter$count = 10004;
	#10 counter$count = 10005;
	#10 counter$count = 10006;
	#10 counter$count = 10007;
	#10 counter$count = 10008;
	#10 counter$count = 10009;
	#10 counter$count = 10010;
	#10 counter$count = 10011;
	#10 counter$count = 10012;
	#10 counter$count = 10013;
	#10 counter$count = 10014;
	#10 counter$count = 10015;
	#10 counter$count = 10016;
	#10 counter$count = 10017;
	#10 counter$count = 10018;
	#10 counter$count = 10019;
	#10 counter$count = 10020;
	#10 counter$count = 10021;
	#10 counter$count = 10022;
	#10 counter$count = 10023;
	#10 counter$count = 10024;
	#10 counter$count = 10025;
	#10 counter$count = 10026;
	#10 counter$count = 10027;
	#10 counter$count = 10028;
	#10 counter$count = 10029;
	#10 counter$count = 10030;
	#10 counter$count = 10031;
	#10 counter$count = 10032;
	#10 counter$count = 10033;
	#10 counter$count = 10034;
	#10 counter$count = 10035;
	#10 counter$count = 10036;
	#10 counter$count = 10037;
	#10 counter$count = 10038;
	#10 counter$count = 10039;
	#10 counter$count = 10040;
	#10 counter$count = 10041;
	#10 counter$count = 10042;
	#10 counter$count = 10043;
	#10 counter$count = 10044;
	#10 counter$count = 10045;
	#10 counter$count = 10046;
	#10 counter$count = 10047;
	#10 counter$count = 10048;
	#10 counter$count = 10049;
	#10 counter$count = 10050;
	#10 counter$count = 10051;
	#10 counter$count = 10052;
	#10 counter$count = 10053;
	#10 counter$count = 10054;
	#10 counter$count = 10055;
	#10 counter$count = 10056;
	#10 counter$count = 10057;
	#10 counter$count = 10058;
	#10 counter$count = 10059;
	#10 counter$count = 10060;
	#10 counter$count = 10061;
	#10 counter$count = 10062;
	#10 counter$count = 10063;
	#10 counter$count = 10064;
	#10 counter$count = 10065;
	#10 counter$count = 10066;
	#10 counter$count = 10067;
	#10 counter$count = 10068;
	#10 counter$count = 10069;
	#10 counter$count = 10070;
	#10 counter$count = 10071;
	#10 counter$count = 10072;
	#10 counter$count = 10073;
	#10 counter$count = 10074;
	#10 counter$count = 10075;
	#10 counter$count = 10076;
	#10 counter$count = 10077;
	#10 counter$count = 10078;
	#10 counter$count = 10079;
	#10 counter$count = 10080;
	#10 counter$count = 10081;
	#10 counter$count = 10082;
	#10 counter$count = 10083;
	#10 counter$count = 10084;
	#10 counter$count = 10085;
	#10 counter$count = 10086;
	#10 counter$count = 10087;
	#10 counter$count = 10088;
	#10 counter$count = 10089;
	#10 counter$count = 10090;
	#10 counter$count = 10091;
	#10 counter$count = 10092;
	#10 counter$count = 10093;
	#10 counter$count = 10094;
	#10 counter$count = 10095;
	#10 counter$count = 10096;
	#10 counter$count = 10097;
	#10 counter$count = 10098;
	#10 counter$count = 10099;
	#10 counter$count = 10100;
	#10 counter$count = 10101;
	#10 counter$count = 10102;
	#10 counter$count = 10103;
	#10 counter$count = 10104;
	#10 counter$count = 10105;
	#10 counter$count = 10106;
	#10 counter$count = 10107;
	#10 counter$count = 10108;
	#10 counter$count = 10109;
	#10 counter$count = 10110;
	#10 counter$count = 10111;
	#10 counter$count = 10112;
	#10 counter$count = 10113;
	#10 counter$count = 10114;
	#10 counter$count = 10115;
	#10 counter$count = 10116;
	#10 counter$count = 10117;
	#10 counter$count = 10118;
	#10 counter$count = 10119;
	#10 counter$count = 10120;
	#10 counter$count = 10121;
	#10 counter$count = 10122;
	#10 counter$count = 10123;
	#10 counter$count = 10124;
	#10 counter$count = 10125;
	#10 counter$count = 10126;
	#10 counter$count = 10127;
	#10 counter$count = 10128;
	#10 counter$count = 10129;
	#10 counter$count = 10130;
	#10 counter$count = 10131;
	#10 counter$count = 10132;
	#10 counter$count = 10133;
	#10 counter$count = 10134;
	#10 counter$count = 10135;
	#10 counter$count = 10136;
	#10 counter$count = 10137;
	#10 counter$count = 10138;
	#10 counter$count = 10139;
	#10 counter$count = 10140;
	#10 counter$count = 10141;
	#10 counter$count = 10142;
	#10 counter$count = 10143;
	#10 counter$count = 10144;
	#10 counter$count = 10145;
	#10 counter$count = 10146;
	#10 counter$count = 10147;
	#10 counter$count = 10148;
	#10 counter$count = 10149;
	#10 counter$count = 10150;
	#10 counter$count = 10151;
	#10 counter$count = 10152;
	#10 counter$count = 10153;
	#10 counter$count = 10154;
	#10 counter$count = 10155;
	#10 counter$count = 10156;
	#10 counter$count = 10157;
	#10 counter$count = 10158;
	#10 counter$count = 10159;
	#10 counter$count = 10160;
	#10 counter$count = 10161;
	#10 counter$count = 10162;
	#10 counter$count = 10163;
	#10 counter$count = 10164;
	#10 counter$count = 10165;
	#10 counter$count = 10166;
	#10 counter$count = 10167;
	#10 counter$count = 10168;
	#10 counter$count = 10169;
	#10 counter$count = 10170;
	#10 counter$count = 10171;
	#10 counter$count = 10172;
	#10 counter$count = 10173;
	#10 counter$count = 10174;
	#10 counter$count = 10175;
	#10 counter$count = 10176;
	#10 counter$count = 10177;
	#10 counter$count = 10178;
	#10 counter$count = 10179;
	#10 counter$count = 10180;
	#10 counter$count = 10181;
	#10 counter$count = 10182;
	#10 counter$count = 10183;
	#10 counter$count = 10184;
	#10 counter$count = 10185;
	#10 counter$count = 10186;
	#10 counter$count = 10187;
	#10 counter$count = 10188;
	#10 counter$count = 10189;
	#10 counter$count = 10190;
	#10 counter$count = 10191;
	#10 counter$count = 10192;
	#10 counter$count = 10193;
	#10 counter$count = 10194;
	#10 counter$count = 10195;
	#10 counter$count = 10196;
	#10 counter$count = 10197;
	#10 counter$count = 10198;
	#10 counter$count = 10199;
	#10 counter$count = 10200;
	#10 counter$count = 10201;
	#10 counter$count = 10202;
	#10 counter$count = 10203;
	#10 counter$count = 10204;
	#10 counter$count = 10205;
	#10 counter$count = 10206;
	#10 counter$count = 10207;
	#10 counter$count = 10208;
	#10 counter$count = 10209;
	#10 counter$count = 10210;
	#10 counter$count = 10211;
	#10 counter$count = 10212;
	#10 counter$count = 10213;
	#10 counter$count = 10214;
	#10 counter$count = 10215;
	#10 counter$count = 10216;
	#10 counter$count = 10217;
	#10 counter$count = 10218;
	#10 counter$count = 10219;
	#10 counter$count = 10220;
	#10 counter$count = 10221;
	#10 counter$count = 10222;
	#10 counter$count = 10223;
	#10 counter$count = 10224;
	#10 counter$count = 10225;
	#10 counter$count = 10226;
	#10 counter$count = 10227;
	#10 counter$count = 10228;
	#10 counter$count = 10229;
	#10 counter$count = 10230;
	#10 counter$count = 10231;
	#10 counter$count = 10232;
	#10 counter$count = 10233;
	#10 counter$count = 10234;
	#10 counter$count = 10235;
	#10 counter$count = 10236;
	#10 counter$count = 10237;
	#10 counter$count = 10238;
	#10 counter$count = 10239;
	#10 counter$count = 10240;
	#10 counter$count = 10241;
	#10 counter$count = 10242;
	#10 counter$count = 10243;
	#10 counter$count = 10244;
	#10 counter$count = 10245;
	#10 counter$count = 10246;
	#10 counter$count = 10247;
	#10 counter$count = 10248;
	#10 counter$count = 10249;
	#10 counter$count = 10250;
	#10 counter$count = 10251;
	#10 counter$count = 10252;
	#10 counter$count = 10253;
	#10 counter$count = 10254;
	#10 counter$count = 10255;
	#10 counter$count = 10256;
	#10 counter$count = 10257;
	#10 counter$count = 10258;
	#10 counter$count = 10259;
	#10 counter$count = 10260;
	#10 counter$count = 10261;
	#10 counter$count = 10262;
	#10 counter$count = 10263;
	#10 counter$count = 10264;
	#10 counter$count = 10265;
	#10 counter$count = 10266;
	#10 counter$count = 10267;
	#10 counter$count = 10268;
	#10 counter$count = 10269;
	#10 counter$count = 10270;
	#10 counter$count = 10271;
	#10 counter$count = 10272;
	#10 counter$count = 10273;
	#10 counter$count = 10274;
	#10 counter$count = 10275;
	#10 counter$count = 10276;
	#10 counter$count = 10277;
	#10 counter$count = 10278;
	#10 counter$count = 10279;
	#10 counter$count = 10280;
	#10 counter$count = 10281;
	#10 counter$count = 10282;
	#10 counter$count = 10283;
	#10 counter$count = 10284;
	#10 counter$count = 10285;
	#10 counter$count = 10286;
	#10 counter$count = 10287;
	#10 counter$count = 10288;
	#10 counter$count = 10289;
	#10 counter$count = 10290;
	#10 counter$count = 10291;
	#10 counter$count = 10292;
	#10 counter$count = 10293;
	#10 counter$count = 10294;
	#10 counter$count = 10295;
	#10 counter$count = 10296;
	#10 counter$count = 10297;
	#10 counter$count = 10298;
	#10 counter$count = 10299;
	#10 counter$count = 10300;
	#10 counter$count = 10301;
	#10 counter$count = 10302;
	#10 counter$count = 10303;
	#10 counter$count = 10304;
	#10 counter$count = 10305;
	#10 counter$count = 10306;
	#10 counter$count = 10307;
	#10 counter$count = 10308;
	#10 counter$count = 10309;
	#10 counter$count = 10310;
	#10 counter$count = 10311;
	#10 counter$count = 10312;
	#10 counter$count = 10313;
	#10 counter$count = 10314;
	#10 counter$count = 10315;
	#10 counter$count = 10316;
	#10 counter$count = 10317;
	#10 counter$count = 10318;
	#10 counter$count = 10319;
	#10 counter$count = 10320;
	#10 counter$count = 10321;
	#10 counter$count = 10322;
	#10 counter$count = 10323;
	#10 counter$count = 10324;
	#10 counter$count = 10325;
	#10 counter$count = 10326;
	#10 counter$count = 10327;
	#10 counter$count = 10328;
	#10 counter$count = 10329;
	#10 counter$count = 10330;
	#10 counter$count = 10331;
	#10 counter$count = 10332;
	#10 counter$count = 10333;
	#10 counter$count = 10334;
	#10 counter$count = 10335;
	#10 counter$count = 10336;
	#10 counter$count = 10337;
	#10 counter$count = 10338;
	#10 counter$count = 10339;
	#10 counter$count = 10340;
	#10 counter$count = 10341;
	#10 counter$count = 10342;
	#10 counter$count = 10343;
	#10 counter$count = 10344;
	#10 counter$count = 10345;
	#10 counter$count = 10346;
	#10 counter$count = 10347;
	#10 counter$count = 10348;
	#10 counter$count = 10349;
	#10 counter$count = 10350;
	#10 counter$count = 10351;
	#10 counter$count = 10352;
	#10 counter$count = 10353;
	#10 counter$count = 10354;
	#10 counter$count = 10355;
	#10 counter$count = 10356;
	#10 counter$count = 10357;
	#10 counter$count = 10358;
	#10 counter$count = 10359;
	#10 counter$count = 10360;
	#10 counter$count = 10361;
	#10 counter$count = 10362;
	#10 counter$count = 10363;
	#10 counter$count = 10364;
	#10 counter$count = 10365;
	#10 counter$count = 10366;
	#10 counter$count = 10367;
	#10 counter$count = 10368;
	#10 counter$count = 10369;
	#10 counter$count = 10370;
	#10 counter$count = 10371;
	#10 counter$count = 10372;
	#10 counter$count = 10373;
	#10 counter$count = 10374;
	#10 counter$count = 10375;
	#10 counter$count = 10376;
	#10 counter$count = 10377;
	#10 counter$count = 10378;
	#10 counter$count = 10379;
	#10 counter$count = 10380;
	#10 counter$count = 10381;
	#10 counter$count = 10382;
	#10 counter$count = 10383;
	#10 counter$count = 10384;
	#10 counter$count = 10385;
	#10 counter$count = 10386;
	#10 counter$count = 10387;
	#10 counter$count = 10388;
	#10 counter$count = 10389;
	#10 counter$count = 10390;
	#10 counter$count = 10391;
	#10 counter$count = 10392;
	#10 counter$count = 10393;
	#10 counter$count = 10394;
	#10 counter$count = 10395;
	#10 counter$count = 10396;
	#10 counter$count = 10397;
	#10 counter$count = 10398;
	#10 counter$count = 10399;
	#10 counter$count = 10400;
	#10 counter$count = 10401;
	#10 counter$count = 10402;
	#10 counter$count = 10403;
	#10 counter$count = 10404;
	#10 counter$count = 10405;
	#10 counter$count = 10406;
	#10 counter$count = 10407;
	#10 counter$count = 10408;
	#10 counter$count = 10409;
	#10 counter$count = 10410;
	#10 counter$count = 10411;
	#10 counter$count = 10412;
	#10 counter$count = 10413;
	#10 counter$count = 10414;
	#10 counter$count = 10415;
	#10 counter$count = 10416;
	#10 counter$count = 10417;
	#10 counter$count = 10418;
	#10 counter$count = 10419;
	#10 counter$count = 10420;
	#10 counter$count = 10421;
	#10 counter$count = 10422;
	#10 counter$count = 10423;
	#10 counter$count = 10424;
	#10 counter$count = 10425;
	#10 counter$count = 10426;
	#10 counter$count = 10427;
	#10 counter$count = 10428;
	#10 counter$count = 10429;
	#10 counter$count = 10430;
	#10 counter$count = 10431;
	#10 counter$count = 10432;
	#10 counter$count = 10433;
	#10 counter$count = 10434;
	#10 counter$count = 10435;
	#10 counter$count = 10436;
	#10 counter$count = 10437;
	#10 counter$count = 10438;
	#10 counter$count = 10439;
	#10 counter$count = 10440;
	#10 counter$count = 10441;
	#10 counter$count = 10442;
	#10 counter$count = 10443;
	#10 counter$count = 10444;
	#10 counter$count = 10445;
	#10 counter$count = 10446;
	#10 counter$count = 10447;
	#10 counter$count = 10448;
	#10 counter$count = 10449;
	#10 counter$count = 10450;
	#10 counter$count = 10451;
	#10 counter$count = 10452;
	#10 counter$count = 10453;
	#10 counter$count = 10454;
	#10 counter$count = 10455;
	#10 counter$count = 10456;
	#10 counter$count = 10457;
	#10 counter$count = 10458;
	#10 counter$count = 10459;
	#10 counter$count = 10460;
	#10 counter$count = 10461;
	#10 counter$count = 10462;
	#10 counter$count = 10463;
	#10 counter$count = 10464;
	#10 counter$count = 10465;
	#10 counter$count = 10466;
	#10 counter$count = 10467;
	#10 counter$count = 10468;
	#10 counter$count = 10469;
	#10 counter$count = 10470;
	#10 counter$count = 10471;
	#10 counter$count = 10472;
	#10 counter$count = 10473;
	#10 counter$count = 10474;
	#10 counter$count = 10475;
	#10 counter$count = 10476;
	#10 counter$count = 10477;
	#10 counter$count = 10478;
	#10 counter$count = 10479;
	#10 counter$count = 10480;
	#10 counter$count = 10481;
	#10 counter$count = 10482;
	#10 counter$count = 10483;
	#10 counter$count = 10484;
	#10 counter$count = 10485;
	#10 counter$count = 10486;
	#10 counter$count = 10487;
	#10 counter$count = 10488;
	#10 counter$count = 10489;
	#10 counter$count = 10490;
	#10 counter$count = 10491;
	#10 counter$count = 10492;
	#10 counter$count = 10493;
	#10 counter$count = 10494;
	#10 counter$count = 10495;
	#10 counter$count = 10496;
	#10 counter$count = 10497;
	#10 counter$count = 10498;
	#10 counter$count = 10499;
	#10 counter$count = 10500;
	#10 counter$count = 10501;
	#10 counter$count = 10502;
	#10 counter$count = 10503;
	#10 counter$count = 10504;
	#10 counter$count = 10505;
	#10 counter$count = 10506;
	#10 counter$count = 10507;
	#10 counter$count = 10508;
	#10 counter$count = 10509;
	#10 counter$count = 10510;
	#10 counter$count = 10511;
	#10 counter$count = 10512;
	#10 counter$count = 10513;
	#10 counter$count = 10514;
	#10 counter$count = 10515;
	#10 counter$count = 10516;
	#10 counter$count = 10517;
	#10 counter$count = 10518;
	#10 counter$count = 10519;
	#10 counter$count = 10520;
	#10 counter$count = 10521;
	#10 counter$count = 10522;
	#10 counter$count = 10523;
	#10 counter$count = 10524;
	#10 counter$count = 10525;
	#10 counter$count = 10526;
	#10 counter$count = 10527;
	#10 counter$count = 10528;
	#10 counter$count = 10529;
	#10 counter$count = 10530;
	#10 counter$count = 10531;
	#10 counter$count = 10532;
	#10 counter$count = 10533;
	#10 counter$count = 10534;
	#10 counter$count = 10535;
	#10 counter$count = 10536;
	#10 counter$count = 10537;
	#10 counter$count = 10538;
	#10 counter$count = 10539;
	#10 counter$count = 10540;
	#10 counter$count = 10541;
	#10 counter$count = 10542;
	#10 counter$count = 10543;
	#10 counter$count = 10544;
	#10 counter$count = 10545;
	#10 counter$count = 10546;
	#10 counter$count = 10547;
	#10 counter$count = 10548;
	#10 counter$count = 10549;
	#10 counter$count = 10550;
	#10 counter$count = 10551;
	#10 counter$count = 10552;
	#10 counter$count = 10553;
	#10 counter$count = 10554;
	#10 counter$count = 10555;
	#10 counter$count = 10556;
	#10 counter$count = 10557;
	#10 counter$count = 10558;
	#10 counter$count = 10559;
	#10 counter$count = 10560;
	#10 counter$count = 10561;
	#10 counter$count = 10562;
	#10 counter$count = 10563;
	#10 counter$count = 10564;
	#10 counter$count = 10565;
	#10 counter$count = 10566;
	#10 counter$count = 10567;
	#10 counter$count = 10568;
	#10 counter$count = 10569;
	#10 counter$count = 10570;
	#10 counter$count = 10571;
	#10 counter$count = 10572;
	#10 counter$count = 10573;
	#10 counter$count = 10574;
	#10 counter$count = 10575;
	#10 counter$count = 10576;
	#10 counter$count = 10577;
	#10 counter$count = 10578;
	#10 counter$count = 10579;
	#10 counter$count = 10580;
	#10 counter$count = 10581;
	#10 counter$count = 10582;
	#10 counter$count = 10583;
	#10 counter$count = 10584;
	#10 counter$count = 10585;
	#10 counter$count = 10586;
	#10 counter$count = 10587;
	#10 counter$count = 10588;
	#10 counter$count = 10589;
	#10 counter$count = 10590;
	#10 counter$count = 10591;
	#10 counter$count = 10592;
	#10 counter$count = 10593;
	#10 counter$count = 10594;
	#10 counter$count = 10595;
	#10 counter$count = 10596;
	#10 counter$count = 10597;
	#10 counter$count = 10598;
	#10 counter$count = 10599;
	#10 counter$count = 10600;
	#10 counter$count = 10601;
	#10 counter$count = 10602;
	#10 counter$count = 10603;
	#10 counter$count = 10604;
	#10 counter$count = 10605;
	#10 counter$count = 10606;
	#10 counter$count = 10607;
	#10 counter$count = 10608;
	#10 counter$count = 10609;
	#10 counter$count = 10610;
	#10 counter$count = 10611;
	#10 counter$count = 10612;
	#10 counter$count = 10613;
	#10 counter$count = 10614;
	#10 counter$count = 10615;
	#10 counter$count = 10616;
	#10 counter$count = 10617;
	#10 counter$count = 10618;
	#10 counter$count = 10619;
	#10 counter$count = 10620;
	#10 counter$count = 10621;
	#10 counter$count = 10622;
	#10 counter$count = 10623;
	#10 counter$count = 10624;
	#10 counter$count = 10625;
	#10 counter$count = 10626;
	#10 counter$count = 10627;
	#10 counter$count = 10628;
	#10 counter$count = 10629;
	#10 counter$count = 10630;
	#10 counter$count = 10631;
	#10 counter$count = 10632;
	#10 counter$count = 10633;
	#10 counter$count = 10634;
	#10 counter$count = 10635;
	#10 counter$count = 10636;
	#10 counter$count = 10637;
	#10 counter$count = 10638;
	#10 counter$count = 10639;
	#10 counter$count = 10640;
	#10 counter$count = 10641;
	#10 counter$count = 10642;
	#10 counter$count = 10643;
	#10 counter$count = 10644;
	#10 counter$count = 10645;
	#10 counter$count = 10646;
	#10 counter$count = 10647;
	#10 counter$count = 10648;
	#10 counter$count = 10649;
	#10 counter$count = 10650;
	#10 counter$count = 10651;
	#10 counter$count = 10652;
	#10 counter$count = 10653;
	#10 counter$count = 10654;
	#10 counter$count = 10655;
	#10 counter$count = 10656;
	#10 counter$count = 10657;
	#10 counter$count = 10658;
	#10 counter$count = 10659;
	#10 counter$count = 10660;
	#10 counter$count = 10661;
	#10 counter$count = 10662;
	#10 counter$count = 10663;
	#10 counter$count = 10664;
	#10 counter$count = 10665;
	#10 counter$count = 10666;
	#10 counter$count = 10667;
	#10 counter$count = 10668;
	#10 counter$count = 10669;
	#10 counter$count = 10670;
	#10 counter$count = 10671;
	#10 counter$count = 10672;
	#10 counter$count = 10673;
	#10 counter$count = 10674;
	#10 counter$count = 10675;
	#10 counter$count = 10676;
	#10 counter$count = 10677;
	#10 counter$count = 10678;
	#10 counter$count = 10679;
	#10 counter$count = 10680;
	#10 counter$count = 10681;
	#10 counter$count = 10682;
	#10 counter$count = 10683;
	#10 counter$count = 10684;
	#10 counter$count = 10685;
	#10 counter$count = 10686;
	#10 counter$count = 10687;
	#10 counter$count = 10688;
	#10 counter$count = 10689;
	#10 counter$count = 10690;
	#10 counter$count = 10691;
	#10 counter$count = 10692;
	#10 counter$count = 10693;
	#10 counter$count = 10694;
	#10 counter$count = 10695;
	#10 counter$count = 10696;
	#10 counter$count = 10697;
	#10 counter$count = 10698;
	#10 counter$count = 10699;
	#10 counter$count = 10700;
	#10 counter$count = 10701;
	#10 counter$count = 10702;
	#10 counter$count = 10703;
	#10 counter$count = 10704;
	#10 counter$count = 10705;
	#10 counter$count = 10706;
	#10 counter$count = 10707;
	#10 counter$count = 10708;
	#10 counter$count = 10709;
	#10 counter$count = 10710;
	#10 counter$count = 10711;
	#10 counter$count = 10712;
	#10 counter$count = 10713;
	#10 counter$count = 10714;
	#10 counter$count = 10715;
	#10 counter$count = 10716;
	#10 counter$count = 10717;
	#10 counter$count = 10718;
	#10 counter$count = 10719;
	#10 counter$count = 10720;
	#10 counter$count = 10721;
	#10 counter$count = 10722;
	#10 counter$count = 10723;
	#10 counter$count = 10724;
	#10 counter$count = 10725;
	#10 counter$count = 10726;
	#10 counter$count = 10727;
	#10 counter$count = 10728;
	#10 counter$count = 10729;
	#10 counter$count = 10730;
	#10 counter$count = 10731;
	#10 counter$count = 10732;
	#10 counter$count = 10733;
	#10 counter$count = 10734;
	#10 counter$count = 10735;
	#10 counter$count = 10736;
	#10 counter$count = 10737;
	#10 counter$count = 10738;
	#10 counter$count = 10739;
	#10 counter$count = 10740;
	#10 counter$count = 10741;
	#10 counter$count = 10742;
	#10 counter$count = 10743;
	#10 counter$count = 10744;
	#10 counter$count = 10745;
	#10 counter$count = 10746;
	#10 counter$count = 10747;
	#10 counter$count = 10748;
	#10 counter$count = 10749;
	#10 counter$count = 10750;
	#10 counter$count = 10751;
	#10 counter$count = 10752;
	#10 counter$count = 10753;
	#10 counter$count = 10754;
	#10 counter$count = 10755;
	#10 counter$count = 10756;
	#10 counter$count = 10757;
	#10 counter$count = 10758;
	#10 counter$count = 10759;
	#10 counter$count = 10760;
	#10 counter$count = 10761;
	#10 counter$count = 10762;
	#10 counter$count = 10763;
	#10 counter$count = 10764;
	#10 counter$count = 10765;
	#10 counter$count = 10766;
	#10 counter$count = 10767;
	#10 counter$count = 10768;
	#10 counter$count = 10769;
	#10 counter$count = 10770;
	#10 counter$count = 10771;
	#10 counter$count = 10772;
	#10 counter$count = 10773;
	#10 counter$count = 10774;
	#10 counter$count = 10775;
	#10 counter$count = 10776;
	#10 counter$count = 10777;
	#10 counter$count = 10778;
	#10 counter$count = 10779;
	#10 counter$count = 10780;
	#10 counter$count = 10781;
	#10 counter$count = 10782;
	#10 counter$count = 10783;
	#10 counter$count = 10784;
	#10 counter$count = 10785;
	#10 counter$count = 10786;
	#10 counter$count = 10787;
	#10 counter$count = 10788;
	#10 counter$count = 10789;
	#10 counter$count = 10790;
	#10 counter$count = 10791;
	#10 counter$count = 10792;
	#10 counter$count = 10793;
	#10 counter$count = 10794;
	#10 counter$count = 10795;
	#10 counter$count = 10796;
	#10 counter$count = 10797;
	#10 counter$count = 10798;
	#10 counter$count = 10799;
	#10 counter$count = 10800;
	#10 counter$count = 10801;
	#10 counter$count = 10802;
	#10 counter$count = 10803;
	#10 counter$count = 10804;
	#10 counter$count = 10805;
	#10 counter$count = 10806;
	#10 counter$count = 10807;
	#10 counter$count = 10808;
	#10 counter$count = 10809;
	#10 counter$count = 10810;
	#10 counter$count = 10811;
	#10 counter$count = 10812;
	#10 counter$count = 10813;
	#10 counter$count = 10814;
	#10 counter$count = 10815;
	#10 counter$count = 10816;
	#10 counter$count = 10817;
	#10 counter$count = 10818;
	#10 counter$count = 10819;
	#10 counter$count = 10820;
	#10 counter$count = 10821;
	#10 counter$count = 10822;
	#10 counter$count = 10823;
	#10 counter$count = 10824;
	#10 counter$count = 10825;
	#10 counter$count = 10826;
	#10 counter$count = 10827;
	#10 counter$count = 10828;
	#10 counter$count = 10829;
	#10 counter$count = 10830;
	#10 counter$count = 10831;
	#10 counter$count = 10832;
	#10 counter$count = 10833;
	#10 counter$count = 10834;
	#10 counter$count = 10835;
	#10 counter$count = 10836;
	#10 counter$count = 10837;
	#10 counter$count = 10838;
	#10 counter$count = 10839;
	#10 counter$count = 10840;
	#10 counter$count = 10841;
	#10 counter$count = 10842;
	#10 counter$count = 10843;
	#10 counter$count = 10844;
	#10 counter$count = 10845;
	#10 counter$count = 10846;
	#10 counter$count = 10847;
	#10 counter$count = 10848;
	#10 counter$count = 10849;
	#10 counter$count = 10850;
	#10 counter$count = 10851;
	#10 counter$count = 10852;
	#10 counter$count = 10853;
	#10 counter$count = 10854;
	#10 counter$count = 10855;
	#10 counter$count = 10856;
	#10 counter$count = 10857;
	#10 counter$count = 10858;
	#10 counter$count = 10859;
	#10 counter$count = 10860;
	#10 counter$count = 10861;
	#10 counter$count = 10862;
	#10 counter$count = 10863;
	#10 counter$count = 10864;
	#10 counter$count = 10865;
	#10 counter$count = 10866;
	#10 counter$count = 10867;
	#10 counter$count = 10868;
	#10 counter$count = 10869;
	#10 counter$count = 10870;
	#10 counter$count = 10871;
	#10 counter$count = 10872;
	#10 counter$count = 10873;
	#10 counter$count = 10874;
	#10 counter$count = 10875;
	#10 counter$count = 10876;
	#10 counter$count = 10877;
	#10 counter$count = 10878;
	#10 counter$count = 10879;
	#10 counter$count = 10880;
	#10 counter$count = 10881;
	#10 counter$count = 10882;
	#10 counter$count = 10883;
	#10 counter$count = 10884;
	#10 counter$count = 10885;
	#10 counter$count = 10886;
	#10 counter$count = 10887;
	#10 counter$count = 10888;
	#10 counter$count = 10889;
	#10 counter$count = 10890;
	#10 counter$count = 10891;
	#10 counter$count = 10892;
	#10 counter$count = 10893;
	#10 counter$count = 10894;
	#10 counter$count = 10895;
	#10 counter$count = 10896;
	#10 counter$count = 10897;
	#10 counter$count = 10898;
	#10 counter$count = 10899;
	#10 counter$count = 10900;
	#10 counter$count = 10901;
	#10 counter$count = 10902;
	#10 counter$count = 10903;
	#10 counter$count = 10904;
	#10 counter$count = 10905;
	#10 counter$count = 10906;
	#10 counter$count = 10907;
	#10 counter$count = 10908;
	#10 counter$count = 10909;
	#10 counter$count = 10910;
	#10 counter$count = 10911;
	#10 counter$count = 10912;
	#10 counter$count = 10913;
	#10 counter$count = 10914;
	#10 counter$count = 10915;
	#10 counter$count = 10916;
	#10 counter$count = 10917;
	#10 counter$count = 10918;
	#10 counter$count = 10919;
	#10 counter$count = 10920;
	#10 counter$count = 10921;
	#10 counter$count = 10922;
	#10 counter$count = 10923;
	#10 counter$count = 10924;
	#10 counter$count = 10925;
	#10 counter$count = 10926;
	#10 counter$count = 10927;
	#10 counter$count = 10928;
	#10 counter$count = 10929;
	#10 counter$count = 10930;
	#10 counter$count = 10931;
	#10 counter$count = 10932;
	#10 counter$count = 10933;
	#10 counter$count = 10934;
	#10 counter$count = 10935;
	#10 counter$count = 10936;
	#10 counter$count = 10937;
	#10 counter$count = 10938;
	#10 counter$count = 10939;
	#10 counter$count = 10940;
	#10 counter$count = 10941;
	#10 counter$count = 10942;
	#10 counter$count = 10943;
	#10 counter$count = 10944;
	#10 counter$count = 10945;
	#10 counter$count = 10946;
	#10 counter$count = 10947;
	#10 counter$count = 10948;
	#10 counter$count = 10949;
	#10 counter$count = 10950;
	#10 counter$count = 10951;
	#10 counter$count = 10952;
	#10 counter$count = 10953;
	#10 counter$count = 10954;
	#10 counter$count = 10955;
	#10 counter$count = 10956;
	#10 counter$count = 10957;
	#10 counter$count = 10958;
	#10 counter$count = 10959;
	#10 counter$count = 10960;
	#10 counter$count = 10961;
	#10 counter$count = 10962;
	#10 counter$count = 10963;
	#10 counter$count = 10964;
	#10 counter$count = 10965;
	#10 counter$count = 10966;
	#10 counter$count = 10967;
	#10 counter$count = 10968;
	#10 counter$count = 10969;
	#10 counter$count = 10970;
	#10 counter$count = 10971;
	#10 counter$count = 10972;
	#10 counter$count = 10973;
	#10 counter$count = 10974;
	#10 counter$count = 10975;
	#10 counter$count = 10976;
	#10 counter$count = 10977;
	#10 counter$count = 10978;
	#10 counter$count = 10979;
	#10 counter$count = 10980;
	#10 counter$count = 10981;
	#10 counter$count = 10982;
	#10 counter$count = 10983;
	#10 counter$count = 10984;
	#10 counter$count = 10985;
	#10 counter$count = 10986;
	#10 counter$count = 10987;
	#10 counter$count = 10988;
	#10 counter$count = 10989;
	#10 counter$count = 10990;
	#10 counter$count = 10991;
	#10 counter$count = 10992;
	#10 counter$count = 10993;
	#10 counter$count = 10994;
	#10 counter$count = 10995;
	#10 counter$count = 10996;
	#10 counter$count = 10997;
	#10 counter$count = 10998;
	#10 counter$count = 10999;
	#10 counter$count = 11000;
	#10 counter$count = 11001;
	#10 counter$count = 11002;
	#10 counter$count = 11003;
	#10 counter$count = 11004;
	#10 counter$count = 11005;
	#10 counter$count = 11006;
	#10 counter$count = 11007;
	#10 counter$count = 11008;
	#10 counter$count = 11009;
	#10 counter$count = 11010;
	#10 counter$count = 11011;
	#10 counter$count = 11012;
	#10 counter$count = 11013;
	#10 counter$count = 11014;
	#10 counter$count = 11015;
	#10 counter$count = 11016;
	#10 counter$count = 11017;
	#10 counter$count = 11018;
	#10 counter$count = 11019;
	#10 counter$count = 11020;
	#10 counter$count = 11021;
	#10 counter$count = 11022;
	#10 counter$count = 11023;
	#10 counter$count = 11024;
	#10 counter$count = 11025;
	#10 counter$count = 11026;
	#10 counter$count = 11027;
	#10 counter$count = 11028;
	#10 counter$count = 11029;
	#10 counter$count = 11030;
	#10 counter$count = 11031;
	#10 counter$count = 11032;
	#10 counter$count = 11033;
	#10 counter$count = 11034;
	#10 counter$count = 11035;
	#10 counter$count = 11036;
	#10 counter$count = 11037;
	#10 counter$count = 11038;
	#10 counter$count = 11039;
	#10 counter$count = 11040;
	#10 counter$count = 11041;
	#10 counter$count = 11042;
	#10 counter$count = 11043;
	#10 counter$count = 11044;
	#10 counter$count = 11045;
	#10 counter$count = 11046;
	#10 counter$count = 11047;
	#10 counter$count = 11048;
	#10 counter$count = 11049;
	#10 counter$count = 11050;
	#10 counter$count = 11051;
	#10 counter$count = 11052;
	#10 counter$count = 11053;
	#10 counter$count = 11054;
	#10 counter$count = 11055;
	#10 counter$count = 11056;
	#10 counter$count = 11057;
	#10 counter$count = 11058;
	#10 counter$count = 11059;
	#10 counter$count = 11060;
	#10 counter$count = 11061;
	#10 counter$count = 11062;
	#10 counter$count = 11063;
	#10 counter$count = 11064;
	#10 counter$count = 11065;
	#10 counter$count = 11066;
	#10 counter$count = 11067;
	#10 counter$count = 11068;
	#10 counter$count = 11069;
	#10 counter$count = 11070;
	#10 counter$count = 11071;
	#10 counter$count = 11072;
	#10 counter$count = 11073;
	#10 counter$count = 11074;
	#10 counter$count = 11075;
	#10 counter$count = 11076;
	#10 counter$count = 11077;
	#10 counter$count = 11078;
	#10 counter$count = 11079;
	#10 counter$count = 11080;
	#10 counter$count = 11081;
	#10 counter$count = 11082;
	#10 counter$count = 11083;
	#10 counter$count = 11084;
	#10 counter$count = 11085;
	#10 counter$count = 11086;
	#10 counter$count = 11087;
	#10 counter$count = 11088;
	#10 counter$count = 11089;
	#10 counter$count = 11090;
	#10 counter$count = 11091;
	#10 counter$count = 11092;
	#10 counter$count = 11093;
	#10 counter$count = 11094;
	#10 counter$count = 11095;
	#10 counter$count = 11096;
	#10 counter$count = 11097;
	#10 counter$count = 11098;
	#10 counter$count = 11099;
	#10 counter$count = 11100;
	#10 counter$count = 11101;
	#10 counter$count = 11102;
	#10 counter$count = 11103;
	#10 counter$count = 11104;
	#10 counter$count = 11105;
	#10 counter$count = 11106;
	#10 counter$count = 11107;
	#10 counter$count = 11108;
	#10 counter$count = 11109;
	#10 counter$count = 11110;
	#10 counter$count = 11111;
	#10 counter$count = 11112;
	#10 counter$count = 11113;
	#10 counter$count = 11114;
	#10 counter$count = 11115;
	#10 counter$count = 11116;
	#10 counter$count = 11117;
	#10 counter$count = 11118;
	#10 counter$count = 11119;
	#10 counter$count = 11120;
	#10 counter$count = 11121;
	#10 counter$count = 11122;
	#10 counter$count = 11123;
	#10 counter$count = 11124;
	#10 counter$count = 11125;
	#10 counter$count = 11126;
	#10 counter$count = 11127;
	#10 counter$count = 11128;
	#10 counter$count = 11129;
	#10 counter$count = 11130;
	#10 counter$count = 11131;
	#10 counter$count = 11132;
	#10 counter$count = 11133;
	#10 counter$count = 11134;
	#10 counter$count = 11135;
	#10 counter$count = 11136;
	#10 counter$count = 11137;
	#10 counter$count = 11138;
	#10 counter$count = 11139;
	#10 counter$count = 11140;
	#10 counter$count = 11141;
	#10 counter$count = 11142;
	#10 counter$count = 11143;
	#10 counter$count = 11144;
	#10 counter$count = 11145;
	#10 counter$count = 11146;
	#10 counter$count = 11147;
	#10 counter$count = 11148;
	#10 counter$count = 11149;
	#10 counter$count = 11150;
	#10 counter$count = 11151;
	#10 counter$count = 11152;
	#10 counter$count = 11153;
	#10 counter$count = 11154;
	#10 counter$count = 11155;
	#10 counter$count = 11156;
	#10 counter$count = 11157;
	#10 counter$count = 11158;
	#10 counter$count = 11159;
	#10 counter$count = 11160;
	#10 counter$count = 11161;
	#10 counter$count = 11162;
	#10 counter$count = 11163;
	#10 counter$count = 11164;
	#10 counter$count = 11165;
	#10 counter$count = 11166;
	#10 counter$count = 11167;
	#10 counter$count = 11168;
	#10 counter$count = 11169;
	#10 counter$count = 11170;
	#10 counter$count = 11171;
	#10 counter$count = 11172;
	#10 counter$count = 11173;
	#10 counter$count = 11174;
	#10 counter$count = 11175;
	#10 counter$count = 11176;
	#10 counter$count = 11177;
	#10 counter$count = 11178;
	#10 counter$count = 11179;
	#10 counter$count = 11180;
	#10 counter$count = 11181;
	#10 counter$count = 11182;
	#10 counter$count = 11183;
	#10 counter$count = 11184;
	#10 counter$count = 11185;
	#10 counter$count = 11186;
	#10 counter$count = 11187;
	#10 counter$count = 11188;
	#10 counter$count = 11189;
	#10 counter$count = 11190;
	#10 counter$count = 11191;
	#10 counter$count = 11192;
	#10 counter$count = 11193;
	#10 counter$count = 11194;
	#10 counter$count = 11195;
	#10 counter$count = 11196;
	#10 counter$count = 11197;
	#10 counter$count = 11198;
	#10 counter$count = 11199;
	#10 counter$count = 11200;
	#10 counter$count = 11201;
	#10 counter$count = 11202;
	#10 counter$count = 11203;
	#10 counter$count = 11204;
	#10 counter$count = 11205;
	#10 counter$count = 11206;
	#10 counter$count = 11207;
	#10 counter$count = 11208;
	#10 counter$count = 11209;
	#10 counter$count = 11210;
	#10 counter$count = 11211;
	#10 counter$count = 11212;
	#10 counter$count = 11213;
	#10 counter$count = 11214;
	#10 counter$count = 11215;
	#10 counter$count = 11216;
	#10 counter$count = 11217;
	#10 counter$count = 11218;
	#10 counter$count = 11219;
	#10 counter$count = 11220;
	#10 counter$count = 11221;
	#10 counter$count = 11222;
	#10 counter$count = 11223;
	#10 counter$count = 11224;
	#10 counter$count = 11225;
	#10 counter$count = 11226;
	#10 counter$count = 11227;
	#10 counter$count = 11228;
	#10 counter$count = 11229;
	#10 counter$count = 11230;
	#10 counter$count = 11231;
	#10 counter$count = 11232;
	#10 counter$count = 11233;
	#10 counter$count = 11234;
	#10 counter$count = 11235;
	#10 counter$count = 11236;
	#10 counter$count = 11237;
	#10 counter$count = 11238;
	#10 counter$count = 11239;
	#10 counter$count = 11240;
	#10 counter$count = 11241;
	#10 counter$count = 11242;
	#10 counter$count = 11243;
	#10 counter$count = 11244;
	#10 counter$count = 11245;
	#10 counter$count = 11246;
	#10 counter$count = 11247;
	#10 counter$count = 11248;
	#10 counter$count = 11249;
	#10 counter$count = 11250;
	#10 counter$count = 11251;
	#10 counter$count = 11252;
	#10 counter$count = 11253;
	#10 counter$count = 11254;
	#10 counter$count = 11255;
	#10 counter$count = 11256;
	#10 counter$count = 11257;
	#10 counter$count = 11258;
	#10 counter$count = 11259;
	#10 counter$count = 11260;
	#10 counter$count = 11261;
	#10 counter$count = 11262;
	#10 counter$count = 11263;
	#10 counter$count = 11264;
	#10 counter$count = 11265;
	#10 counter$count = 11266;
	#10 counter$count = 11267;
	#10 counter$count = 11268;
	#10 counter$count = 11269;
	#10 counter$count = 11270;
	#10 counter$count = 11271;
	#10 counter$count = 11272;
	#10 counter$count = 11273;
	#10 counter$count = 11274;
	#10 counter$count = 11275;
	#10 counter$count = 11276;
	#10 counter$count = 11277;
	#10 counter$count = 11278;
	#10 counter$count = 11279;
	#10 counter$count = 11280;
	#10 counter$count = 11281;
	#10 counter$count = 11282;
	#10 counter$count = 11283;
	#10 counter$count = 11284;
	#10 counter$count = 11285;
	#10 counter$count = 11286;
	#10 counter$count = 11287;
	#10 counter$count = 11288;
	#10 counter$count = 11289;
	#10 counter$count = 11290;
	#10 counter$count = 11291;
	#10 counter$count = 11292;
	#10 counter$count = 11293;
	#10 counter$count = 11294;
	#10 counter$count = 11295;
	#10 counter$count = 11296;
	#10 counter$count = 11297;
	#10 counter$count = 11298;
	#10 counter$count = 11299;
	#10 counter$count = 11300;
	#10 counter$count = 11301;
	#10 counter$count = 11302;
	#10 counter$count = 11303;
	#10 counter$count = 11304;
	#10 counter$count = 11305;
	#10 counter$count = 11306;
	#10 counter$count = 11307;
	#10 counter$count = 11308;
	#10 counter$count = 11309;
	#10 counter$count = 11310;
	#10 counter$count = 11311;
	#10 counter$count = 11312;
	#10 counter$count = 11313;
	#10 counter$count = 11314;
	#10 counter$count = 11315;
	#10 counter$count = 11316;
	#10 counter$count = 11317;
	#10 counter$count = 11318;
	#10 counter$count = 11319;
	#10 counter$count = 11320;
	#10 counter$count = 11321;
	#10 counter$count = 11322;
	#10 counter$count = 11323;
	#10 counter$count = 11324;
	#10 counter$count = 11325;
	#10 counter$count = 11326;
	#10 counter$count = 11327;
	#10 counter$count = 11328;
	#10 counter$count = 11329;
	#10 counter$count = 11330;
	#10 counter$count = 11331;
	#10 counter$count = 11332;
	#10 counter$count = 11333;
	#10 counter$count = 11334;
	#10 counter$count = 11335;
	#10 counter$count = 11336;
	#10 counter$count = 11337;
	#10 counter$count = 11338;
	#10 counter$count = 11339;
	#10 counter$count = 11340;
	#10 counter$count = 11341;
	#10 counter$count = 11342;
	#10 counter$count = 11343;
	#10 counter$count = 11344;
	#10 counter$count = 11345;
	#10 counter$count = 11346;
	#10 counter$count = 11347;
	#10 counter$count = 11348;
	#10 counter$count = 11349;
	#10 counter$count = 11350;
	#10 counter$count = 11351;
	#10 counter$count = 11352;
	#10 counter$count = 11353;
	#10 counter$count = 11354;
	#10 counter$count = 11355;
	#10 counter$count = 11356;
	#10 counter$count = 11357;
	#10 counter$count = 11358;
	#10 counter$count = 11359;
	#10 counter$count = 11360;
	#10 counter$count = 11361;
	#10 counter$count = 11362;
	#10 counter$count = 11363;
	#10 counter$count = 11364;
	#10 counter$count = 11365;
	#10 counter$count = 11366;
	#10 counter$count = 11367;
	#10 counter$count = 11368;
	#10 counter$count = 11369;
	#10 counter$count = 11370;
	#10 counter$count = 11371;
	#10 counter$count = 11372;
	#10 counter$count = 11373;
	#10 counter$count = 11374;
	#10 counter$count = 11375;
	#10 counter$count = 11376;
	#10 counter$count = 11377;
	#10 counter$count = 11378;
	#10 counter$count = 11379;
	#10 counter$count = 11380;
	#10 counter$count = 11381;
	#10 counter$count = 11382;
	#10 counter$count = 11383;
	#10 counter$count = 11384;
	#10 counter$count = 11385;
	#10 counter$count = 11386;
	#10 counter$count = 11387;
	#10 counter$count = 11388;
	#10 counter$count = 11389;
	#10 counter$count = 11390;
	#10 counter$count = 11391;
	#10 counter$count = 11392;
	#10 counter$count = 11393;
	#10 counter$count = 11394;
	#10 counter$count = 11395;
	#10 counter$count = 11396;
	#10 counter$count = 11397;
	#10 counter$count = 11398;
	#10 counter$count = 11399;
	#10 counter$count = 11400;
	#10 counter$count = 11401;
	#10 counter$count = 11402;
	#10 counter$count = 11403;
	#10 counter$count = 11404;
	#10 counter$count = 11405;
	#10 counter$count = 11406;
	#10 counter$count = 11407;
	#10 counter$count = 11408;
	#10 counter$count = 11409;
	#10 counter$count = 11410;
	#10 counter$count = 11411;
	#10 counter$count = 11412;
	#10 counter$count = 11413;
	#10 counter$count = 11414;
	#10 counter$count = 11415;
	#10 counter$count = 11416;
	#10 counter$count = 11417;
	#10 counter$count = 11418;
	#10 counter$count = 11419;
	#10 counter$count = 11420;
	#10 counter$count = 11421;
	#10 counter$count = 11422;
	#10 counter$count = 11423;
	#10 counter$count = 11424;
	#10 counter$count = 11425;
	#10 counter$count = 11426;
	#10 counter$count = 11427;
	#10 counter$count = 11428;
	#10 counter$count = 11429;
	#10 counter$count = 11430;
	#10 counter$count = 11431;
	#10 counter$count = 11432;
	#10 counter$count = 11433;
	#10 counter$count = 11434;
	#10 counter$count = 11435;
	#10 counter$count = 11436;
	#10 counter$count = 11437;
	#10 counter$count = 11438;
	#10 counter$count = 11439;
	#10 counter$count = 11440;
	#10 counter$count = 11441;
	#10 counter$count = 11442;
	#10 counter$count = 11443;
	#10 counter$count = 11444;
	#10 counter$count = 11445;
	#10 counter$count = 11446;
	#10 counter$count = 11447;
	#10 counter$count = 11448;
	#10 counter$count = 11449;
	#10 counter$count = 11450;
	#10 counter$count = 11451;
	#10 counter$count = 11452;
	#10 counter$count = 11453;
	#10 counter$count = 11454;
	#10 counter$count = 11455;
	#10 counter$count = 11456;
	#10 counter$count = 11457;
	#10 counter$count = 11458;
	#10 counter$count = 11459;
	#10 counter$count = 11460;
	#10 counter$count = 11461;
	#10 counter$count = 11462;
	#10 counter$count = 11463;
	#10 counter$count = 11464;
	#10 counter$count = 11465;
	#10 counter$count = 11466;
	#10 counter$count = 11467;
	#10 counter$count = 11468;
	#10 counter$count = 11469;
	#10 counter$count = 11470;
	#10 counter$count = 11471;
	#10 counter$count = 11472;
	#10 counter$count = 11473;
	#10 counter$count = 11474;
	#10 counter$count = 11475;
	#10 counter$count = 11476;
	#10 counter$count = 11477;
	#10 counter$count = 11478;
	#10 counter$count = 11479;
	#10 counter$count = 11480;
	#10 counter$count = 11481;
	#10 counter$count = 11482;
	#10 counter$count = 11483;
	#10 counter$count = 11484;
	#10 counter$count = 11485;
	#10 counter$count = 11486;
	#10 counter$count = 11487;
	#10 counter$count = 11488;
	#10 counter$count = 11489;
	#10 counter$count = 11490;
	#10 counter$count = 11491;
	#10 counter$count = 11492;
	#10 counter$count = 11493;
	#10 counter$count = 11494;
	#10 counter$count = 11495;
	#10 counter$count = 11496;
	#10 counter$count = 11497;
	#10 counter$count = 11498;
	#10 counter$count = 11499;
	#10 counter$count = 11500;
	#10 counter$count = 11501;
	#10 counter$count = 11502;
	#10 counter$count = 11503;
	#10 counter$count = 11504;
	#10 counter$count = 11505;
	#10 counter$count = 11506;
	#10 counter$count = 11507;
	#10 counter$count = 11508;
	#10 counter$count = 11509;
	#10 counter$count = 11510;
	#10 counter$count = 11511;
	#10 counter$count = 11512;
	#10 counter$count = 11513;
	#10 counter$count = 11514;
	#10 counter$count = 11515;
	#10 counter$count = 11516;
	#10 counter$count = 11517;
	#10 counter$count = 11518;
	#10 counter$count = 11519;
	#10 counter$count = 11520;
	#10 counter$count = 11521;
	#10 counter$count = 11522;
	#10 counter$count = 11523;
	#10 counter$count = 11524;
	#10 counter$count = 11525;
	#10 counter$count = 11526;
	#10 counter$count = 11527;
	#10 counter$count = 11528;
	#10 counter$count = 11529;
	#10 counter$count = 11530;
	#10 counter$count = 11531;
	#10 counter$count = 11532;
	#10 counter$count = 11533;
	#10 counter$count = 11534;
	#10 counter$count = 11535;
	#10 counter$count = 11536;
	#10 counter$count = 11537;
	#10 counter$count = 11538;
	#10 counter$count = 11539;
	#10 counter$count = 11540;
	#10 counter$count = 11541;
	#10 counter$count = 11542;
	#10 counter$count = 11543;
	#10 counter$count = 11544;
	#10 counter$count = 11545;
	#10 counter$count = 11546;
	#10 counter$count = 11547;
	#10 counter$count = 11548;
	#10 counter$count = 11549;
	#10 counter$count = 11550;
	#10 counter$count = 11551;
	#10 counter$count = 11552;
	#10 counter$count = 11553;
	#10 counter$count = 11554;
	#10 counter$count = 11555;
	#10 counter$count = 11556;
	#10 counter$count = 11557;
	#10 counter$count = 11558;
	#10 counter$count = 11559;
	#10 counter$count = 11560;
	#10 counter$count = 11561;
	#10 counter$count = 11562;
	#10 counter$count = 11563;
	#10 counter$count = 11564;
	#10 counter$count = 11565;
	#10 counter$count = 11566;
	#10 counter$count = 11567;
	#10 counter$count = 11568;
	#10 counter$count = 11569;
	#10 counter$count = 11570;
	#10 counter$count = 11571;
	#10 counter$count = 11572;
	#10 counter$count = 11573;
	#10 counter$count = 11574;
	#10 counter$count = 11575;
	#10 counter$count = 11576;
	#10 counter$count = 11577;
	#10 counter$count = 11578;
	#10 counter$count = 11579;
	#10 counter$count = 11580;
	#10 counter$count = 11581;
	#10 counter$count = 11582;
	#10 counter$count = 11583;
	#10 counter$count = 11584;
	#10 counter$count = 11585;
	#10 counter$count = 11586;
	#10 counter$count = 11587;
	#10 counter$count = 11588;
	#10 counter$count = 11589;
	#10 counter$count = 11590;
	#10 counter$count = 11591;
	#10 counter$count = 11592;
	#10 counter$count = 11593;
	#10 counter$count = 11594;
	#10 counter$count = 11595;
	#10 counter$count = 11596;
	#10 counter$count = 11597;
	#10 counter$count = 11598;
	#10 counter$count = 11599;
	#10 counter$count = 11600;
	#10 counter$count = 11601;
	#10 counter$count = 11602;
	#10 counter$count = 11603;
	#10 counter$count = 11604;
	#10 counter$count = 11605;
	#10 counter$count = 11606;
	#10 counter$count = 11607;
	#10 counter$count = 11608;
	#10 counter$count = 11609;
	#10 counter$count = 11610;
	#10 counter$count = 11611;
	#10 counter$count = 11612;
	#10 counter$count = 11613;
	#10 counter$count = 11614;
	#10 counter$count = 11615;
	#10 counter$count = 11616;
	#10 counter$count = 11617;
	#10 counter$count = 11618;
	#10 counter$count = 11619;
	#10 counter$count = 11620;
	#10 counter$count = 11621;
	#10 counter$count = 11622;
	#10 counter$count = 11623;
	#10 counter$count = 11624;
	#10 counter$count = 11625;
	#10 counter$count = 11626;
	#10 counter$count = 11627;
	#10 counter$count = 11628;
	#10 counter$count = 11629;
	#10 counter$count = 11630;
	#10 counter$count = 11631;
	#10 counter$count = 11632;
	#10 counter$count = 11633;
	#10 counter$count = 11634;
	#10 counter$count = 11635;
	#10 counter$count = 11636;
	#10 counter$count = 11637;
	#10 counter$count = 11638;
	#10 counter$count = 11639;
	#10 counter$count = 11640;
	#10 counter$count = 11641;
	#10 counter$count = 11642;
	#10 counter$count = 11643;
	#10 counter$count = 11644;
	#10 counter$count = 11645;
	#10 counter$count = 11646;
	#10 counter$count = 11647;
	#10 counter$count = 11648;
	#10 counter$count = 11649;
	#10 counter$count = 11650;
	#10 counter$count = 11651;
	#10 counter$count = 11652;
	#10 counter$count = 11653;
	#10 counter$count = 11654;
	#10 counter$count = 11655;
	#10 counter$count = 11656;
	#10 counter$count = 11657;
	#10 counter$count = 11658;
	#10 counter$count = 11659;
	#10 counter$count = 11660;
	#10 counter$count = 11661;
	#10 counter$count = 11662;
	#10 counter$count = 11663;
	#10 counter$count = 11664;
	#10 counter$count = 11665;
	#10 counter$count = 11666;
	#10 counter$count = 11667;
	#10 counter$count = 11668;
	#10 counter$count = 11669;
	#10 counter$count = 11670;
	#10 counter$count = 11671;
	#10 counter$count = 11672;
	#10 counter$count = 11673;
	#10 counter$count = 11674;
	#10 counter$count = 11675;
	#10 counter$count = 11676;
	#10 counter$count = 11677;
	#10 counter$count = 11678;
	#10 counter$count = 11679;
	#10 counter$count = 11680;
	#10 counter$count = 11681;
	#10 counter$count = 11682;
	#10 counter$count = 11683;
	#10 counter$count = 11684;
	#10 counter$count = 11685;
	#10 counter$count = 11686;
	#10 counter$count = 11687;
	#10 counter$count = 11688;
	#10 counter$count = 11689;
	#10 counter$count = 11690;
	#10 counter$count = 11691;
	#10 counter$count = 11692;
	#10 counter$count = 11693;
	#10 counter$count = 11694;
	#10 counter$count = 11695;
	#10 counter$count = 11696;
	#10 counter$count = 11697;
	#10 counter$count = 11698;
	#10 counter$count = 11699;
	#10 counter$count = 11700;
	#10 counter$count = 11701;
	#10 counter$count = 11702;
	#10 counter$count = 11703;
	#10 counter$count = 11704;
	#10 counter$count = 11705;
	#10 counter$count = 11706;
	#10 counter$count = 11707;
	#10 counter$count = 11708;
	#10 counter$count = 11709;
	#10 counter$count = 11710;
	#10 counter$count = 11711;
	#10 counter$count = 11712;
	#10 counter$count = 11713;
	#10 counter$count = 11714;
	#10 counter$count = 11715;
	#10 counter$count = 11716;
	#10 counter$count = 11717;
	#10 counter$count = 11718;
	#10 counter$count = 11719;
	#10 counter$count = 11720;
	#10 counter$count = 11721;
	#10 counter$count = 11722;
	#10 counter$count = 11723;
	#10 counter$count = 11724;
	#10 counter$count = 11725;
	#10 counter$count = 11726;
	#10 counter$count = 11727;
	#10 counter$count = 11728;
	#10 counter$count = 11729;
	#10 counter$count = 11730;
	#10 counter$count = 11731;
	#10 counter$count = 11732;
	#10 counter$count = 11733;
	#10 counter$count = 11734;
	#10 counter$count = 11735;
	#10 counter$count = 11736;
	#10 counter$count = 11737;
	#10 counter$count = 11738;
	#10 counter$count = 11739;
	#10 counter$count = 11740;
	#10 counter$count = 11741;
	#10 counter$count = 11742;
	#10 counter$count = 11743;
	#10 counter$count = 11744;
	#10 counter$count = 11745;
	#10 counter$count = 11746;
	#10 counter$count = 11747;
	#10 counter$count = 11748;
	#10 counter$count = 11749;
	#10 counter$count = 11750;
	#10 counter$count = 11751;
	#10 counter$count = 11752;
	#10 counter$count = 11753;
	#10 counter$count = 11754;
	#10 counter$count = 11755;
	#10 counter$count = 11756;
	#10 counter$count = 11757;
	#10 counter$count = 11758;
	#10 counter$count = 11759;
	#10 counter$count = 11760;
	#10 counter$count = 11761;
	#10 counter$count = 11762;
	#10 counter$count = 11763;
	#10 counter$count = 11764;
	#10 counter$count = 11765;
	#10 counter$count = 11766;
	#10 counter$count = 11767;
	#10 counter$count = 11768;
	#10 counter$count = 11769;
	#10 counter$count = 11770;
	#10 counter$count = 11771;
	#10 counter$count = 11772;
	#10 counter$count = 11773;
	#10 counter$count = 11774;
	#10 counter$count = 11775;
	#10 counter$count = 11776;
	#10 counter$count = 11777;
	#10 counter$count = 11778;
	#10 counter$count = 11779;
	#10 counter$count = 11780;
	#10 counter$count = 11781;
	#10 counter$count = 11782;
	#10 counter$count = 11783;
	#10 counter$count = 11784;
	#10 counter$count = 11785;
	#10 counter$count = 11786;
	#10 counter$count = 11787;
	#10 counter$count = 11788;
	#10 counter$count = 11789;
	#10 counter$count = 11790;
	#10 counter$count = 11791;
	#10 counter$count = 11792;
	#10 counter$count = 11793;
	#10 counter$count = 11794;
	#10 counter$count = 11795;
	#10 counter$count = 11796;
	#10 counter$count = 11797;
	#10 counter$count = 11798;
	#10 counter$count = 11799;
	#10 counter$count = 11800;
	#10 counter$count = 11801;
	#10 counter$count = 11802;
	#10 counter$count = 11803;
	#10 counter$count = 11804;
	#10 counter$count = 11805;
	#10 counter$count = 11806;
	#10 counter$count = 11807;
	#10 counter$count = 11808;
	#10 counter$count = 11809;
	#10 counter$count = 11810;
	#10 counter$count = 11811;
	#10 counter$count = 11812;
	#10 counter$count = 11813;
	#10 counter$count = 11814;
	#10 counter$count = 11815;
	#10 counter$count = 11816;
	#10 counter$count = 11817;
	#10 counter$count = 11818;
	#10 counter$count = 11819;
	#10 counter$count = 11820;
	#10 counter$count = 11821;
	#10 counter$count = 11822;
	#10 counter$count = 11823;
	#10 counter$count = 11824;
	#10 counter$count = 11825;
	#10 counter$count = 11826;
	#10 counter$count = 11827;
	#10 counter$count = 11828;
	#10 counter$count = 11829;
	#10 counter$count = 11830;
	#10 counter$count = 11831;
	#10 counter$count = 11832;
	#10 counter$count = 11833;
	#10 counter$count = 11834;
	#10 counter$count = 11835;
	#10 counter$count = 11836;
	#10 counter$count = 11837;
	#10 counter$count = 11838;
	#10 counter$count = 11839;
	#10 counter$count = 11840;
	#10 counter$count = 11841;
	#10 counter$count = 11842;
	#10 counter$count = 11843;
	#10 counter$count = 11844;
	#10 counter$count = 11845;
	#10 counter$count = 11846;
	#10 counter$count = 11847;
	#10 counter$count = 11848;
	#10 counter$count = 11849;
	#10 counter$count = 11850;
	#10 counter$count = 11851;
	#10 counter$count = 11852;
	#10 counter$count = 11853;
	#10 counter$count = 11854;
	#10 counter$count = 11855;
	#10 counter$count = 11856;
	#10 counter$count = 11857;
	#10 counter$count = 11858;
	#10 counter$count = 11859;
	#10 counter$count = 11860;
	#10 counter$count = 11861;
	#10 counter$count = 11862;
	#10 counter$count = 11863;
	#10 counter$count = 11864;
	#10 counter$count = 11865;
	#10 counter$count = 11866;
	#10 counter$count = 11867;
	#10 counter$count = 11868;
	#10 counter$count = 11869;
	#10 counter$count = 11870;
	#10 counter$count = 11871;
	#10 counter$count = 11872;
	#10 counter$count = 11873;
	#10 counter$count = 11874;
	#10 counter$count = 11875;
	#10 counter$count = 11876;
	#10 counter$count = 11877;
	#10 counter$count = 11878;
	#10 counter$count = 11879;
	#10 counter$count = 11880;
	#10 counter$count = 11881;
	#10 counter$count = 11882;
	#10 counter$count = 11883;
	#10 counter$count = 11884;
	#10 counter$count = 11885;
	#10 counter$count = 11886;
	#10 counter$count = 11887;
	#10 counter$count = 11888;
	#10 counter$count = 11889;
	#10 counter$count = 11890;
	#10 counter$count = 11891;
	#10 counter$count = 11892;
	#10 counter$count = 11893;
	#10 counter$count = 11894;
	#10 counter$count = 11895;
	#10 counter$count = 11896;
	#10 counter$count = 11897;
	#10 counter$count = 11898;
	#10 counter$count = 11899;
	#10 counter$count = 11900;
	#10 counter$count = 11901;
	#10 counter$count = 11902;
	#10 counter$count = 11903;
	#10 counter$count = 11904;
	#10 counter$count = 11905;
	#10 counter$count = 11906;
	#10 counter$count = 11907;
	#10 counter$count = 11908;
	#10 counter$count = 11909;
	#10 counter$count = 11910;
	#10 counter$count = 11911;
	#10 counter$count = 11912;
	#10 counter$count = 11913;
	#10 counter$count = 11914;
	#10 counter$count = 11915;
	#10 counter$count = 11916;
	#10 counter$count = 11917;
	#10 counter$count = 11918;
	#10 counter$count = 11919;
	#10 counter$count = 11920;
	#10 counter$count = 11921;
	#10 counter$count = 11922;
	#10 counter$count = 11923;
	#10 counter$count = 11924;
	#10 counter$count = 11925;
	#10 counter$count = 11926;
	#10 counter$count = 11927;
	#10 counter$count = 11928;
	#10 counter$count = 11929;
	#10 counter$count = 11930;
	#10 counter$count = 11931;
	#10 counter$count = 11932;
	#10 counter$count = 11933;
	#10 counter$count = 11934;
	#10 counter$count = 11935;
	#10 counter$count = 11936;
	#10 counter$count = 11937;
	#10 counter$count = 11938;
	#10 counter$count = 11939;
	#10 counter$count = 11940;
	#10 counter$count = 11941;
	#10 counter$count = 11942;
	#10 counter$count = 11943;
	#10 counter$count = 11944;
	#10 counter$count = 11945;
	#10 counter$count = 11946;
	#10 counter$count = 11947;
	#10 counter$count = 11948;
	#10 counter$count = 11949;
	#10 counter$count = 11950;
	#10 counter$count = 11951;
	#10 counter$count = 11952;
	#10 counter$count = 11953;
	#10 counter$count = 11954;
	#10 counter$count = 11955;
	#10 counter$count = 11956;
	#10 counter$count = 11957;
	#10 counter$count = 11958;
	#10 counter$count = 11959;
	#10 counter$count = 11960;
	#10 counter$count = 11961;
	#10 counter$count = 11962;
	#10 counter$count = 11963;
	#10 counter$count = 11964;
	#10 counter$count = 11965;
	#10 counter$count = 11966;
	#10 counter$count = 11967;
	#10 counter$count = 11968;
	#10 counter$count = 11969;
	#10 counter$count = 11970;
	#10 counter$count = 11971;
	#10 counter$count = 11972;
	#10 counter$count = 11973;
	#10 counter$count = 11974;
	#10 counter$count = 11975;
	#10 counter$count = 11976;
	#10 counter$count = 11977;
	#10 counter$count = 11978;
	#10 counter$count = 11979;
	#10 counter$count = 11980;
	#10 counter$count = 11981;
	#10 counter$count = 11982;
	#10 counter$count = 11983;
	#10 counter$count = 11984;
	#10 counter$count = 11985;
	#10 counter$count = 11986;
	#10 counter$count = 11987;
	#10 counter$count = 11988;
	#10 counter$count = 11989;
	#10 counter$count = 11990;
	#10 counter$count = 11991;
	#10 counter$count = 11992;
	#10 counter$count = 11993;
	#10 counter$count = 11994;
	#10 counter$count = 11995;
	#10 counter$count = 11996;
	#10 counter$count = 11997;
	#10 counter$count = 11998;
	#10 counter$count = 11999;
	#10 counter$count = 12000;
	#10 counter$count = 12001;
	#10 counter$count = 12002;
	#10 counter$count = 12003;
	#10 counter$count = 12004;
	#10 counter$count = 12005;
	#10 counter$count = 12006;
	#10 counter$count = 12007;
	#10 counter$count = 12008;
	#10 counter$count = 12009;
	#10 counter$count = 12010;
	#10 counter$count = 12011;
	#10 counter$count = 12012;
	#10 counter$count = 12013;
	#10 counter$count = 12014;
	#10 counter$count = 12015;
	#10 counter$count = 12016;
	#10 counter$count = 12017;
	#10 counter$count = 12018;
	#10 counter$count = 12019;
	#10 counter$count = 12020;
	#10 counter$count = 12021;
	#10 counter$count = 12022;
	#10 counter$count = 12023;
	#10 counter$count = 12024;
	#10 counter$count = 12025;
	#10 counter$count = 12026;
	#10 counter$count = 12027;
	#10 counter$count = 12028;
	#10 counter$count = 12029;
	#10 counter$count = 12030;
	#10 counter$count = 12031;
	#10 counter$count = 12032;
	#10 counter$count = 12033;
	#10 counter$count = 12034;
	#10 counter$count = 12035;
	#10 counter$count = 12036;
	#10 counter$count = 12037;
	#10 counter$count = 12038;
	#10 counter$count = 12039;
	#10 counter$count = 12040;
	#10 counter$count = 12041;
	#10 counter$count = 12042;
	#10 counter$count = 12043;
	#10 counter$count = 12044;
	#10 counter$count = 12045;
	#10 counter$count = 12046;
	#10 counter$count = 12047;
	#10 counter$count = 12048;
	#10 counter$count = 12049;
	#10 counter$count = 12050;
	#10 counter$count = 12051;
	#10 counter$count = 12052;
	#10 counter$count = 12053;
	#10 counter$count = 12054;
	#10 counter$count = 12055;
	#10 counter$count = 12056;
	#10 counter$count = 12057;
	#10 counter$count = 12058;
	#10 counter$count = 12059;
	#10 counter$count = 12060;
	#10 counter$count = 12061;
	#10 counter$count = 12062;
	#10 counter$count = 12063;
	#10 counter$count = 12064;
	#10 counter$count = 12065;
	#10 counter$count = 12066;
	#10 counter$count = 12067;
	#10 counter$count = 12068;
	#10 counter$count = 12069;
	#10 counter$count = 12070;
	#10 counter$count = 12071;
	#10 counter$count = 12072;
	#10 counter$count = 12073;
	#10 counter$count = 12074;
	#10 counter$count = 12075;
	#10 counter$count = 12076;
	#10 counter$count = 12077;
	#10 counter$count = 12078;
	#10 counter$count = 12079;
	#10 counter$count = 12080;
	#10 counter$count = 12081;
	#10 counter$count = 12082;
	#10 counter$count = 12083;
	#10 counter$count = 12084;
	#10 counter$count = 12085;
	#10 counter$count = 12086;
	#10 counter$count = 12087;
	#10 counter$count = 12088;
	#10 counter$count = 12089;
	#10 counter$count = 12090;
	#10 counter$count = 12091;
	#10 counter$count = 12092;
	#10 counter$count = 12093;
	#10 counter$count = 12094;
	#10 counter$count = 12095;
	#10 counter$count = 12096;
	#10 counter$count = 12097;
	#10 counter$count = 12098;
	#10 counter$count = 12099;
	#10 counter$count = 12100;
	#10 counter$count = 12101;
	#10 counter$count = 12102;
	#10 counter$count = 12103;
	#10 counter$count = 12104;
	#10 counter$count = 12105;
	#10 counter$count = 12106;
	#10 counter$count = 12107;
	#10 counter$count = 12108;
	#10 counter$count = 12109;
	#10 counter$count = 12110;
	#10 counter$count = 12111;
	#10 counter$count = 12112;
	#10 counter$count = 12113;
	#10 counter$count = 12114;
	#10 counter$count = 12115;
	#10 counter$count = 12116;
	#10 counter$count = 12117;
	#10 counter$count = 12118;
	#10 counter$count = 12119;
	#10 counter$count = 12120;
	#10 counter$count = 12121;
	#10 counter$count = 12122;
	#10 counter$count = 12123;
	#10 counter$count = 12124;
	#10 counter$count = 12125;
	#10 counter$count = 12126;
	#10 counter$count = 12127;
	#10 counter$count = 12128;
	#10 counter$count = 12129;
	#10 counter$count = 12130;
	#10 counter$count = 12131;
	#10 counter$count = 12132;
	#10 counter$count = 12133;
	#10 counter$count = 12134;
	#10 counter$count = 12135;
	#10 counter$count = 12136;
	#10 counter$count = 12137;
	#10 counter$count = 12138;
	#10 counter$count = 12139;
	#10 counter$count = 12140;
	#10 counter$count = 12141;
	#10 counter$count = 12142;
	#10 counter$count = 12143;
	#10 counter$count = 12144;
	#10 counter$count = 12145;
	#10 counter$count = 12146;
	#10 counter$count = 12147;
	#10 counter$count = 12148;
	#10 counter$count = 12149;
	#10 counter$count = 12150;
	#10 counter$count = 12151;
	#10 counter$count = 12152;
	#10 counter$count = 12153;
	#10 counter$count = 12154;
	#10 counter$count = 12155;
	#10 counter$count = 12156;
	#10 counter$count = 12157;
	#10 counter$count = 12158;
	#10 counter$count = 12159;
	#10 counter$count = 12160;
	#10 counter$count = 12161;
	#10 counter$count = 12162;
	#10 counter$count = 12163;
	#10 counter$count = 12164;
	#10 counter$count = 12165;
	#10 counter$count = 12166;
	#10 counter$count = 12167;
	#10 counter$count = 12168;
	#10 counter$count = 12169;
	#10 counter$count = 12170;
	#10 counter$count = 12171;
	#10 counter$count = 12172;
	#10 counter$count = 12173;
	#10 counter$count = 12174;
	#10 counter$count = 12175;
	#10 counter$count = 12176;
	#10 counter$count = 12177;
	#10 counter$count = 12178;
	#10 counter$count = 12179;
	#10 counter$count = 12180;
	#10 counter$count = 12181;
	#10 counter$count = 12182;
	#10 counter$count = 12183;
	#10 counter$count = 12184;
	#10 counter$count = 12185;
	#10 counter$count = 12186;
	#10 counter$count = 12187;
	#10 counter$count = 12188;
	#10 counter$count = 12189;
	#10 counter$count = 12190;
	#10 counter$count = 12191;
	#10 counter$count = 12192;
	#10 counter$count = 12193;
	#10 counter$count = 12194;
	#10 counter$count = 12195;
	#10 counter$count = 12196;
	#10 counter$count = 12197;
	#10 counter$count = 12198;
	#10 counter$count = 12199;
	#10 counter$count = 12200;
	#10 counter$count = 12201;
	#10 counter$count = 12202;
	#10 counter$count = 12203;
	#10 counter$count = 12204;
	#10 counter$count = 12205;
	#10 counter$count = 12206;
	#10 counter$count = 12207;
	#10 counter$count = 12208;
	#10 counter$count = 12209;
	#10 counter$count = 12210;
	#10 counter$count = 12211;
	#10 counter$count = 12212;
	#10 counter$count = 12213;
	#10 counter$count = 12214;
	#10 counter$count = 12215;
	#10 counter$count = 12216;
	#10 counter$count = 12217;
	#10 counter$count = 12218;
	#10 counter$count = 12219;
	#10 counter$count = 12220;
	#10 counter$count = 12221;
	#10 counter$count = 12222;
	#10 counter$count = 12223;
	#10 counter$count = 12224;
	#10 counter$count = 12225;
	#10 counter$count = 12226;
	#10 counter$count = 12227;
	#10 counter$count = 12228;
	#10 counter$count = 12229;
	#10 counter$count = 12230;
	#10 counter$count = 12231;
	#10 counter$count = 12232;
	#10 counter$count = 12233;
	#10 counter$count = 12234;
	#10 counter$count = 12235;
	#10 counter$count = 12236;
	#10 counter$count = 12237;
	#10 counter$count = 12238;
	#10 counter$count = 12239;
	#10 counter$count = 12240;
	#10 counter$count = 12241;
	#10 counter$count = 12242;
	#10 counter$count = 12243;
	#10 counter$count = 12244;
	#10 counter$count = 12245;
	#10 counter$count = 12246;
	#10 counter$count = 12247;
	#10 counter$count = 12248;
	#10 counter$count = 12249;
	#10 counter$count = 12250;
	#10 counter$count = 12251;
	#10 counter$count = 12252;
	#10 counter$count = 12253;
	#10 counter$count = 12254;
	#10 counter$count = 12255;
	#10 counter$count = 12256;
	#10 counter$count = 12257;
	#10 counter$count = 12258;
	#10 counter$count = 12259;
	#10 counter$count = 12260;
	#10 counter$count = 12261;
	#10 counter$count = 12262;
	#10 counter$count = 12263;
	#10 counter$count = 12264;
	#10 counter$count = 12265;
	#10 counter$count = 12266;
	#10 counter$count = 12267;
	#10 counter$count = 12268;
	#10 counter$count = 12269;
	#10 counter$count = 12270;
	#10 counter$count = 12271;
	#10 counter$count = 12272;
	#10 counter$count = 12273;
	#10 counter$count = 12274;
	#10 counter$count = 12275;
	#10 counter$count = 12276;
	#10 counter$count = 12277;
	#10 counter$count = 12278;
	#10 counter$count = 12279;
	#10 counter$count = 12280;
	#10 counter$count = 12281;
	#10 counter$count = 12282;
	#10 counter$count = 12283;
	#10 counter$count = 12284;
	#10 counter$count = 12285;
	#10 counter$count = 12286;
	#10 counter$count = 12287;
	#10 counter$count = 12288;
	#10 counter$count = 12289;
	#10 counter$count = 12290;
	#10 counter$count = 12291;
	#10 counter$count = 12292;
	#10 counter$count = 12293;
	#10 counter$count = 12294;
	#10 counter$count = 12295;
	#10 counter$count = 12296;
	#10 counter$count = 12297;
	#10 counter$count = 12298;
	#10 counter$count = 12299;
	#10 counter$count = 12300;
	#10 counter$count = 12301;
	#10 counter$count = 12302;
	#10 counter$count = 12303;
	#10 counter$count = 12304;
	#10 counter$count = 12305;
	#10 counter$count = 12306;
	#10 counter$count = 12307;
	#10 counter$count = 12308;
	#10 counter$count = 12309;
	#10 counter$count = 12310;
	#10 counter$count = 12311;
	#10 counter$count = 12312;
	#10 counter$count = 12313;
	#10 counter$count = 12314;
	#10 counter$count = 12315;
	#10 counter$count = 12316;
	#10 counter$count = 12317;
	#10 counter$count = 12318;
	#10 counter$count = 12319;
	#10 counter$count = 12320;
	#10 counter$count = 12321;
	#10 counter$count = 12322;
	#10 counter$count = 12323;
	#10 counter$count = 12324;
	#10 counter$count = 12325;
	#10 counter$count = 12326;
	#10 counter$count = 12327;
	#10 counter$count = 12328;
	#10 counter$count = 12329;
	#10 counter$count = 12330;
	#10 counter$count = 12331;
	#10 counter$count = 12332;
	#10 counter$count = 12333;
	#10 counter$count = 12334;
	#10 counter$count = 12335;
	#10 counter$count = 12336;
	#10 counter$count = 12337;
	#10 counter$count = 12338;
	#10 counter$count = 12339;
	#10 counter$count = 12340;
	#10 counter$count = 12341;
	#10 counter$count = 12342;
	#10 counter$count = 12343;
	#10 counter$count = 12344;
	#10 counter$count = 12345;
	#10 counter$count = 12346;
	#10 counter$count = 12347;
	#10 counter$count = 12348;
	#10 counter$count = 12349;
	#10 counter$count = 12350;
	#10 counter$count = 12351;
	#10 counter$count = 12352;
	#10 counter$count = 12353;
	#10 counter$count = 12354;
	#10 counter$count = 12355;
	#10 counter$count = 12356;
	#10 counter$count = 12357;
	#10 counter$count = 12358;
	#10 counter$count = 12359;
	#10 counter$count = 12360;
	#10 counter$count = 12361;
	#10 counter$count = 12362;
	#10 counter$count = 12363;
	#10 counter$count = 12364;
	#10 counter$count = 12365;
	#10 counter$count = 12366;
	#10 counter$count = 12367;
	#10 counter$count = 12368;
	#10 counter$count = 12369;
	#10 counter$count = 12370;
	#10 counter$count = 12371;
	#10 counter$count = 12372;
	#10 counter$count = 12373;
	#10 counter$count = 12374;
	#10 counter$count = 12375;
	#10 counter$count = 12376;
	#10 counter$count = 12377;
	#10 counter$count = 12378;
	#10 counter$count = 12379;
	#10 counter$count = 12380;
	#10 counter$count = 12381;
	#10 counter$count = 12382;
	#10 counter$count = 12383;
	#10 counter$count = 12384;
	#10 counter$count = 12385;
	#10 counter$count = 12386;
	#10 counter$count = 12387;
	#10 counter$count = 12388;
	#10 counter$count = 12389;
	#10 counter$count = 12390;
	#10 counter$count = 12391;
	#10 counter$count = 12392;
	#10 counter$count = 12393;
	#10 counter$count = 12394;
	#10 counter$count = 12395;
	#10 counter$count = 12396;
	#10 counter$count = 12397;
	#10 counter$count = 12398;
	#10 counter$count = 12399;
	#10 counter$count = 12400;
	#10 counter$count = 12401;
	#10 counter$count = 12402;
	#10 counter$count = 12403;
	#10 counter$count = 12404;
	#10 counter$count = 12405;
	#10 counter$count = 12406;
	#10 counter$count = 12407;
	#10 counter$count = 12408;
	#10 counter$count = 12409;
	#10 counter$count = 12410;
	#10 counter$count = 12411;
	#10 counter$count = 12412;
	#10 counter$count = 12413;
	#10 counter$count = 12414;
	#10 counter$count = 12415;
	#10 counter$count = 12416;
	#10 counter$count = 12417;
	#10 counter$count = 12418;
	#10 counter$count = 12419;
	#10 counter$count = 12420;
	#10 counter$count = 12421;
	#10 counter$count = 12422;
	#10 counter$count = 12423;
	#10 counter$count = 12424;
	#10 counter$count = 12425;
	#10 counter$count = 12426;
	#10 counter$count = 12427;
	#10 counter$count = 12428;
	#10 counter$count = 12429;
	#10 counter$count = 12430;
	#10 counter$count = 12431;
	#10 counter$count = 12432;
	#10 counter$count = 12433;
	#10 counter$count = 12434;
	#10 counter$count = 12435;
	#10 counter$count = 12436;
	#10 counter$count = 12437;
	#10 counter$count = 12438;
	#10 counter$count = 12439;
	#10 counter$count = 12440;
	#10 counter$count = 12441;
	#10 counter$count = 12442;
	#10 counter$count = 12443;
	#10 counter$count = 12444;
	#10 counter$count = 12445;
	#10 counter$count = 12446;
	#10 counter$count = 12447;
	#10 counter$count = 12448;
	#10 counter$count = 12449;
	#10 counter$count = 12450;
	#10 counter$count = 12451;
	#10 counter$count = 12452;
	#10 counter$count = 12453;
	#10 counter$count = 12454;
	#10 counter$count = 12455;
	#10 counter$count = 12456;
	#10 counter$count = 12457;
	#10 counter$count = 12458;
	#10 counter$count = 12459;
	#10 counter$count = 12460;
	#10 counter$count = 12461;
	#10 counter$count = 12462;
	#10 counter$count = 12463;
	#10 counter$count = 12464;
	#10 counter$count = 12465;
	#10 counter$count = 12466;
	#10 counter$count = 12467;
	#10 counter$count = 12468;
	#10 counter$count = 12469;
	#10 counter$count = 12470;
	#10 counter$count = 12471;
	#10 counter$count = 12472;
	#10 counter$count = 12473;
	#10 counter$count = 12474;
	#10 counter$count = 12475;
	#10 counter$count = 12476;
	#10 counter$count = 12477;
	#10 counter$count = 12478;
	#10 counter$count = 12479;
	#10 counter$count = 12480;
	#10 counter$count = 12481;
	#10 counter$count = 12482;
	#10 counter$count = 12483;
	#10 counter$count = 12484;
	#10 counter$count = 12485;
	#10 counter$count = 12486;
	#10 counter$count = 12487;
	#10 counter$count = 12488;
	#10 counter$count = 12489;
	#10 counter$count = 12490;
	#10 counter$count = 12491;
	#10 counter$count = 12492;
	#10 counter$count = 12493;
	#10 counter$count = 12494;
	#10 counter$count = 12495;
	#10 counter$count = 12496;
	#10 counter$count = 12497;
	#10 counter$count = 12498;
	#10 counter$count = 12499;
	#10 counter$count = 12500;
	#10 counter$count = 12501;
	#10 counter$count = 12502;
	#10 counter$count = 12503;
	#10 counter$count = 12504;
	#10 counter$count = 12505;
	#10 counter$count = 12506;
	#10 counter$count = 12507;
	#10 counter$count = 12508;
	#10 counter$count = 12509;
	#10 counter$count = 12510;
	#10 counter$count = 12511;
	#10 counter$count = 12512;
	#10 counter$count = 12513;
	#10 counter$count = 12514;
	#10 counter$count = 12515;
	#10 counter$count = 12516;
	#10 counter$count = 12517;
	#10 counter$count = 12518;
	#10 counter$count = 12519;
	#10 counter$count = 12520;
	#10 counter$count = 12521;
	#10 counter$count = 12522;
	#10 counter$count = 12523;
	#10 counter$count = 12524;
	#10 counter$count = 12525;
	#10 counter$count = 12526;
	#10 counter$count = 12527;
	#10 counter$count = 12528;
	#10 counter$count = 12529;
	#10 counter$count = 12530;
	#10 counter$count = 12531;
	#10 counter$count = 12532;
	#10 counter$count = 12533;
	#10 counter$count = 12534;
	#10 counter$count = 12535;
	#10 counter$count = 12536;
	#10 counter$count = 12537;
	#10 counter$count = 12538;
	#10 counter$count = 12539;
	#10 counter$count = 12540;
	#10 counter$count = 12541;
	#10 counter$count = 12542;
	#10 counter$count = 12543;
	#10 counter$count = 12544;
	#10 counter$count = 12545;
	#10 counter$count = 12546;
	#10 counter$count = 12547;
	#10 counter$count = 12548;
	#10 counter$count = 12549;
	#10 counter$count = 12550;
	#10 counter$count = 12551;
	#10 counter$count = 12552;
	#10 counter$count = 12553;
	#10 counter$count = 12554;
	#10 counter$count = 12555;
	#10 counter$count = 12556;
	#10 counter$count = 12557;
	#10 counter$count = 12558;
	#10 counter$count = 12559;
	#10 counter$count = 12560;
	#10 counter$count = 12561;
	#10 counter$count = 12562;
	#10 counter$count = 12563;
	#10 counter$count = 12564;
	#10 counter$count = 12565;
	#10 counter$count = 12566;
	#10 counter$count = 12567;
	#10 counter$count = 12568;
	#10 counter$count = 12569;
	#10 counter$count = 12570;
	#10 counter$count = 12571;
	#10 counter$count = 12572;
	#10 counter$count = 12573;
	#10 counter$count = 12574;
	#10 counter$count = 12575;
	#10 counter$count = 12576;
	#10 counter$count = 12577;
	#10 counter$count = 12578;
	#10 counter$count = 12579;
	#10 counter$count = 12580;
	#10 counter$count = 12581;
	#10 counter$count = 12582;
	#10 counter$count = 12583;
	#10 counter$count = 12584;
	#10 counter$count = 12585;
	#10 counter$count = 12586;
	#10 counter$count = 12587;
	#10 counter$count = 12588;
	#10 counter$count = 12589;
	#10 counter$count = 12590;
	#10 counter$count = 12591;
	#10 counter$count = 12592;
	#10 counter$count = 12593;
	#10 counter$count = 12594;
	#10 counter$count = 12595;
	#10 counter$count = 12596;
	#10 counter$count = 12597;
	#10 counter$count = 12598;
	#10 counter$count = 12599;
	#10 counter$count = 12600;
	#10 counter$count = 12601;
	#10 counter$count = 12602;
	#10 counter$count = 12603;
	#10 counter$count = 12604;
	#10 counter$count = 12605;
	#10 counter$count = 12606;
	#10 counter$count = 12607;
	#10 counter$count = 12608;
	#10 counter$count = 12609;
	#10 counter$count = 12610;
	#10 counter$count = 12611;
	#10 counter$count = 12612;
	#10 counter$count = 12613;
	#10 counter$count = 12614;
	#10 counter$count = 12615;
	#10 counter$count = 12616;
	#10 counter$count = 12617;
	#10 counter$count = 12618;
	#10 counter$count = 12619;
	#10 counter$count = 12620;
	#10 counter$count = 12621;
	#10 counter$count = 12622;
	#10 counter$count = 12623;
	#10 counter$count = 12624;
	#10 counter$count = 12625;
	#10 counter$count = 12626;
	#10 counter$count = 12627;
	#10 counter$count = 12628;
	#10 counter$count = 12629;
	#10 counter$count = 12630;
	#10 counter$count = 12631;
	#10 counter$count = 12632;
	#10 counter$count = 12633;
	#10 counter$count = 12634;
	#10 counter$count = 12635;
	#10 counter$count = 12636;
	#10 counter$count = 12637;
	#10 counter$count = 12638;
	#10 counter$count = 12639;
	#10 counter$count = 12640;
	#10 counter$count = 12641;
	#10 counter$count = 12642;
	#10 counter$count = 12643;
	#10 counter$count = 12644;
	#10 counter$count = 12645;
	#10 counter$count = 12646;
	#10 counter$count = 12647;
	#10 counter$count = 12648;
	#10 counter$count = 12649;
	#10 counter$count = 12650;
	#10 counter$count = 12651;
	#10 counter$count = 12652;
	#10 counter$count = 12653;
	#10 counter$count = 12654;
	#10 counter$count = 12655;
	#10 counter$count = 12656;
	#10 counter$count = 12657;
	#10 counter$count = 12658;
	#10 counter$count = 12659;
	#10 counter$count = 12660;
	#10 counter$count = 12661;
	#10 counter$count = 12662;
	#10 counter$count = 12663;
	#10 counter$count = 12664;
	#10 counter$count = 12665;
	#10 counter$count = 12666;
	#10 counter$count = 12667;
	#10 counter$count = 12668;
	#10 counter$count = 12669;
	#10 counter$count = 12670;
	#10 counter$count = 12671;
	#10 counter$count = 12672;
	#10 counter$count = 12673;
	#10 counter$count = 12674;
	#10 counter$count = 12675;
	#10 counter$count = 12676;
	#10 counter$count = 12677;
	#10 counter$count = 12678;
	#10 counter$count = 12679;
	#10 counter$count = 12680;
	#10 counter$count = 12681;
	#10 counter$count = 12682;
	#10 counter$count = 12683;
	#10 counter$count = 12684;
	#10 counter$count = 12685;
	#10 counter$count = 12686;
	#10 counter$count = 12687;
	#10 counter$count = 12688;
	#10 counter$count = 12689;
	#10 counter$count = 12690;
	#10 counter$count = 12691;
	#10 counter$count = 12692;
	#10 counter$count = 12693;
	#10 counter$count = 12694;
	#10 counter$count = 12695;
	#10 counter$count = 12696;
	#10 counter$count = 12697;
	#10 counter$count = 12698;
	#10 counter$count = 12699;
	#10 counter$count = 12700;
	#10 counter$count = 12701;
	#10 counter$count = 12702;
	#10 counter$count = 12703;
	#10 counter$count = 12704;
	#10 counter$count = 12705;
	#10 counter$count = 12706;
	#10 counter$count = 12707;
	#10 counter$count = 12708;
	#10 counter$count = 12709;
	#10 counter$count = 12710;
	#10 counter$count = 12711;
	#10 counter$count = 12712;
	#10 counter$count = 12713;
	#10 counter$count = 12714;
	#10 counter$count = 12715;
	#10 counter$count = 12716;
	#10 counter$count = 12717;
	#10 counter$count = 12718;
	#10 counter$count = 12719;
	#10 counter$count = 12720;
	#10 counter$count = 12721;
	#10 counter$count = 12722;
	#10 counter$count = 12723;
	#10 counter$count = 12724;
	#10 counter$count = 12725;
	#10 counter$count = 12726;
	#10 counter$count = 12727;
	#10 counter$count = 12728;
	#10 counter$count = 12729;
	#10 counter$count = 12730;
	#10 counter$count = 12731;
	#10 counter$count = 12732;
	#10 counter$count = 12733;
	#10 counter$count = 12734;
	#10 counter$count = 12735;
	#10 counter$count = 12736;
	#10 counter$count = 12737;
	#10 counter$count = 12738;
	#10 counter$count = 12739;
	#10 counter$count = 12740;
	#10 counter$count = 12741;
	#10 counter$count = 12742;
	#10 counter$count = 12743;
	#10 counter$count = 12744;
	#10 counter$count = 12745;
	#10 counter$count = 12746;
	#10 counter$count = 12747;
	#10 counter$count = 12748;
	#10 counter$count = 12749;
	#10 counter$count = 12750;
	#10 counter$count = 12751;
	#10 counter$count = 12752;
	#10 counter$count = 12753;
	#10 counter$count = 12754;
	#10 counter$count = 12755;
	#10 counter$count = 12756;
	#10 counter$count = 12757;
	#10 counter$count = 12758;
	#10 counter$count = 12759;
	#10 counter$count = 12760;
	#10 counter$count = 12761;
	#10 counter$count = 12762;
	#10 counter$count = 12763;
	#10 counter$count = 12764;
	#10 counter$count = 12765;
	#10 counter$count = 12766;
	#10 counter$count = 12767;
	#10 counter$count = 12768;
	#10 counter$count = 12769;
	#10 counter$count = 12770;
	#10 counter$count = 12771;
	#10 counter$count = 12772;
	#10 counter$count = 12773;
	#10 counter$count = 12774;
	#10 counter$count = 12775;
	#10 counter$count = 12776;
	#10 counter$count = 12777;
	#10 counter$count = 12778;
	#10 counter$count = 12779;
	#10 counter$count = 12780;
	#10 counter$count = 12781;
	#10 counter$count = 12782;
	#10 counter$count = 12783;
	#10 counter$count = 12784;
	#10 counter$count = 12785;
	#10 counter$count = 12786;
	#10 counter$count = 12787;
	#10 counter$count = 12788;
	#10 counter$count = 12789;
	#10 counter$count = 12790;
	#10 counter$count = 12791;
	#10 counter$count = 12792;
	#10 counter$count = 12793;
	#10 counter$count = 12794;
	#10 counter$count = 12795;
	#10 counter$count = 12796;
	#10 counter$count = 12797;
	#10 counter$count = 12798;
	#10 counter$count = 12799;
	#10 counter$count = 12800;
	#10 counter$count = 12801;
	#10 counter$count = 12802;
	#10 counter$count = 12803;
	#10 counter$count = 12804;
	#10 counter$count = 12805;
	#10 counter$count = 12806;
	#10 counter$count = 12807;
	#10 counter$count = 12808;
	#10 counter$count = 12809;
	#10 counter$count = 12810;
	#10 counter$count = 12811;
	#10 counter$count = 12812;
	#10 counter$count = 12813;
	#10 counter$count = 12814;
	#10 counter$count = 12815;
	#10 counter$count = 12816;
	#10 counter$count = 12817;
	#10 counter$count = 12818;
	#10 counter$count = 12819;
	#10 counter$count = 12820;
	#10 counter$count = 12821;
	#10 counter$count = 12822;
	#10 counter$count = 12823;
	#10 counter$count = 12824;
	#10 counter$count = 12825;
	#10 counter$count = 12826;
	#10 counter$count = 12827;
	#10 counter$count = 12828;
	#10 counter$count = 12829;
	#10 counter$count = 12830;
	#10 counter$count = 12831;
	#10 counter$count = 12832;
	#10 counter$count = 12833;
	#10 counter$count = 12834;
	#10 counter$count = 12835;
	#10 counter$count = 12836;
	#10 counter$count = 12837;
	#10 counter$count = 12838;
	#10 counter$count = 12839;
	#10 counter$count = 12840;
	#10 counter$count = 12841;
	#10 counter$count = 12842;
	#10 counter$count = 12843;
	#10 counter$count = 12844;
	#10 counter$count = 12845;
	#10 counter$count = 12846;
	#10 counter$count = 12847;
	#10 counter$count = 12848;
	#10 counter$count = 12849;
	#10 counter$count = 12850;
	#10 counter$count = 12851;
	#10 counter$count = 12852;
	#10 counter$count = 12853;
	#10 counter$count = 12854;
	#10 counter$count = 12855;
	#10 counter$count = 12856;
	#10 counter$count = 12857;
	#10 counter$count = 12858;
	#10 counter$count = 12859;
	#10 counter$count = 12860;
	#10 counter$count = 12861;
	#10 counter$count = 12862;
	#10 counter$count = 12863;
	#10 counter$count = 12864;
	#10 counter$count = 12865;
	#10 counter$count = 12866;
	#10 counter$count = 12867;
	#10 counter$count = 12868;
	#10 counter$count = 12869;
	#10 counter$count = 12870;
	#10 counter$count = 12871;
	#10 counter$count = 12872;
	#10 counter$count = 12873;
	#10 counter$count = 12874;
	#10 counter$count = 12875;
	#10 counter$count = 12876;
	#10 counter$count = 12877;
	#10 counter$count = 12878;
	#10 counter$count = 12879;
	#10 counter$count = 12880;
	#10 counter$count = 12881;
	#10 counter$count = 12882;
	#10 counter$count = 12883;
	#10 counter$count = 12884;
	#10 counter$count = 12885;
	#10 counter$count = 12886;
	#10 counter$count = 12887;
	#10 counter$count = 12888;
	#10 counter$count = 12889;
	#10 counter$count = 12890;
	#10 counter$count = 12891;
	#10 counter$count = 12892;
	#10 counter$count = 12893;
	#10 counter$count = 12894;
	#10 counter$count = 12895;
	#10 counter$count = 12896;
	#10 counter$count = 12897;
	#10 counter$count = 12898;
	#10 counter$count = 12899;
	#10 counter$count = 12900;
	#10 counter$count = 12901;
	#10 counter$count = 12902;
	#10 counter$count = 12903;
	#10 counter$count = 12904;
	#10 counter$count = 12905;
	#10 counter$count = 12906;
	#10 counter$count = 12907;
	#10 counter$count = 12908;
	#10 counter$count = 12909;
	#10 counter$count = 12910;
	#10 counter$count = 12911;
	#10 counter$count = 12912;
	#10 counter$count = 12913;
	#10 counter$count = 12914;
	#10 counter$count = 12915;
	#10 counter$count = 12916;
	#10 counter$count = 12917;
	#10 counter$count = 12918;
	#10 counter$count = 12919;
	#10 counter$count = 12920;
	#10 counter$count = 12921;
	#10 counter$count = 12922;
	#10 counter$count = 12923;
	#10 counter$count = 12924;
	#10 counter$count = 12925;
	#10 counter$count = 12926;
	#10 counter$count = 12927;
	#10 counter$count = 12928;
	#10 counter$count = 12929;
	#10 counter$count = 12930;
	#10 counter$count = 12931;
	#10 counter$count = 12932;
	#10 counter$count = 12933;
	#10 counter$count = 12934;
	#10 counter$count = 12935;
	#10 counter$count = 12936;
	#10 counter$count = 12937;
	#10 counter$count = 12938;
	#10 counter$count = 12939;
	#10 counter$count = 12940;
	#10 counter$count = 12941;
	#10 counter$count = 12942;
	#10 counter$count = 12943;
	#10 counter$count = 12944;
	#10 counter$count = 12945;
	#10 counter$count = 12946;
	#10 counter$count = 12947;
	#10 counter$count = 12948;
	#10 counter$count = 12949;
	#10 counter$count = 12950;
	#10 counter$count = 12951;
	#10 counter$count = 12952;
	#10 counter$count = 12953;
	#10 counter$count = 12954;
	#10 counter$count = 12955;
	#10 counter$count = 12956;
	#10 counter$count = 12957;
	#10 counter$count = 12958;
	#10 counter$count = 12959;
	#10 counter$count = 12960;
	#10 counter$count = 12961;
	#10 counter$count = 12962;
	#10 counter$count = 12963;
	#10 counter$count = 12964;
	#10 counter$count = 12965;
	#10 counter$count = 12966;
	#10 counter$count = 12967;
	#10 counter$count = 12968;
	#10 counter$count = 12969;
	#10 counter$count = 12970;
	#10 counter$count = 12971;
	#10 counter$count = 12972;
	#10 counter$count = 12973;
	#10 counter$count = 12974;
	#10 counter$count = 12975;
	#10 counter$count = 12976;
	#10 counter$count = 12977;
	#10 counter$count = 12978;
	#10 counter$count = 12979;
	#10 counter$count = 12980;
	#10 counter$count = 12981;
	#10 counter$count = 12982;
	#10 counter$count = 12983;
	#10 counter$count = 12984;
	#10 counter$count = 12985;
	#10 counter$count = 12986;
	#10 counter$count = 12987;
	#10 counter$count = 12988;
	#10 counter$count = 12989;
	#10 counter$count = 12990;
	#10 counter$count = 12991;
	#10 counter$count = 12992;
	#10 counter$count = 12993;
	#10 counter$count = 12994;
	#10 counter$count = 12995;
	#10 counter$count = 12996;
	#10 counter$count = 12997;
	#10 counter$count = 12998;
	#10 counter$count = 12999;
	#10 counter$count = 13000;
	#10 counter$count = 13001;
	#10 counter$count = 13002;
	#10 counter$count = 13003;
	#10 counter$count = 13004;
	#10 counter$count = 13005;
	#10 counter$count = 13006;
	#10 counter$count = 13007;
	#10 counter$count = 13008;
	#10 counter$count = 13009;
	#10 counter$count = 13010;
	#10 counter$count = 13011;
	#10 counter$count = 13012;
	#10 counter$count = 13013;
	#10 counter$count = 13014;
	#10 counter$count = 13015;
	#10 counter$count = 13016;
	#10 counter$count = 13017;
	#10 counter$count = 13018;
	#10 counter$count = 13019;
	#10 counter$count = 13020;
	#10 counter$count = 13021;
	#10 counter$count = 13022;
	#10 counter$count = 13023;
	#10 counter$count = 13024;
	#10 counter$count = 13025;
	#10 counter$count = 13026;
	#10 counter$count = 13027;
	#10 counter$count = 13028;
	#10 counter$count = 13029;
	#10 counter$count = 13030;
	#10 counter$count = 13031;
	#10 counter$count = 13032;
	#10 counter$count = 13033;
	#10 counter$count = 13034;
	#10 counter$count = 13035;
	#10 counter$count = 13036;
	#10 counter$count = 13037;
	#10 counter$count = 13038;
	#10 counter$count = 13039;
	#10 counter$count = 13040;
	#10 counter$count = 13041;
	#10 counter$count = 13042;
	#10 counter$count = 13043;
	#10 counter$count = 13044;
	#10 counter$count = 13045;
	#10 counter$count = 13046;
	#10 counter$count = 13047;
	#10 counter$count = 13048;
	#10 counter$count = 13049;
	#10 counter$count = 13050;
	#10 counter$count = 13051;
	#10 counter$count = 13052;
	#10 counter$count = 13053;
	#10 counter$count = 13054;
	#10 counter$count = 13055;
	#10 counter$count = 13056;
	#10 counter$count = 13057;
	#10 counter$count = 13058;
	#10 counter$count = 13059;
	#10 counter$count = 13060;
	#10 counter$count = 13061;
	#10 counter$count = 13062;
	#10 counter$count = 13063;
	#10 counter$count = 13064;
	#10 counter$count = 13065;
	#10 counter$count = 13066;
	#10 counter$count = 13067;
	#10 counter$count = 13068;
	#10 counter$count = 13069;
	#10 counter$count = 13070;
	#10 counter$count = 13071;
	#10 counter$count = 13072;
	#10 counter$count = 13073;
	#10 counter$count = 13074;
	#10 counter$count = 13075;
	#10 counter$count = 13076;
	#10 counter$count = 13077;
	#10 counter$count = 13078;
	#10 counter$count = 13079;
	#10 counter$count = 13080;
	#10 counter$count = 13081;
	#10 counter$count = 13082;
	#10 counter$count = 13083;
	#10 counter$count = 13084;
	#10 counter$count = 13085;
	#10 counter$count = 13086;
	#10 counter$count = 13087;
	#10 counter$count = 13088;
	#10 counter$count = 13089;
	#10 counter$count = 13090;
	#10 counter$count = 13091;
	#10 counter$count = 13092;
	#10 counter$count = 13093;
	#10 counter$count = 13094;
	#10 counter$count = 13095;
	#10 counter$count = 13096;
	#10 counter$count = 13097;
	#10 counter$count = 13098;
	#10 counter$count = 13099;
	#10 counter$count = 13100;
	#10 counter$count = 13101;
	#10 counter$count = 13102;
	#10 counter$count = 13103;
	#10 counter$count = 13104;
	#10 counter$count = 13105;
	#10 counter$count = 13106;
	#10 counter$count = 13107;
	#10 counter$count = 13108;
	#10 counter$count = 13109;
	#10 counter$count = 13110;
	#10 counter$count = 13111;
	#10 counter$count = 13112;
	#10 counter$count = 13113;
	#10 counter$count = 13114;
	#10 counter$count = 13115;
	#10 counter$count = 13116;
	#10 counter$count = 13117;
	#10 counter$count = 13118;
	#10 counter$count = 13119;
	#10 counter$count = 13120;
	#10 counter$count = 13121;
	#10 counter$count = 13122;
	#10 counter$count = 13123;
	#10 counter$count = 13124;
	#10 counter$count = 13125;
	#10 counter$count = 13126;
	#10 counter$count = 13127;
	#10 counter$count = 13128;
	#10 counter$count = 13129;
	#10 counter$count = 13130;
	#10 counter$count = 13131;
	#10 counter$count = 13132;
	#10 counter$count = 13133;
	#10 counter$count = 13134;
	#10 counter$count = 13135;
	#10 counter$count = 13136;
	#10 counter$count = 13137;
	#10 counter$count = 13138;
	#10 counter$count = 13139;
	#10 counter$count = 13140;
	#10 counter$count = 13141;
	#10 counter$count = 13142;
	#10 counter$count = 13143;
	#10 counter$count = 13144;
	#10 counter$count = 13145;
	#10 counter$count = 13146;
	#10 counter$count = 13147;
	#10 counter$count = 13148;
	#10 counter$count = 13149;
	#10 counter$count = 13150;
	#10 counter$count = 13151;
	#10 counter$count = 13152;
	#10 counter$count = 13153;
	#10 counter$count = 13154;
	#10 counter$count = 13155;
	#10 counter$count = 13156;
	#10 counter$count = 13157;
	#10 counter$count = 13158;
	#10 counter$count = 13159;
	#10 counter$count = 13160;
	#10 counter$count = 13161;
	#10 counter$count = 13162;
	#10 counter$count = 13163;
	#10 counter$count = 13164;
	#10 counter$count = 13165;
	#10 counter$count = 13166;
	#10 counter$count = 13167;
	#10 counter$count = 13168;
	#10 counter$count = 13169;
	#10 counter$count = 13170;
	#10 counter$count = 13171;
	#10 counter$count = 13172;
	#10 counter$count = 13173;
	#10 counter$count = 13174;
	#10 counter$count = 13175;
	#10 counter$count = 13176;
	#10 counter$count = 13177;
	#10 counter$count = 13178;
	#10 counter$count = 13179;
	#10 counter$count = 13180;
	#10 counter$count = 13181;
	#10 counter$count = 13182;
	#10 counter$count = 13183;
	#10 counter$count = 13184;
	#10 counter$count = 13185;
	#10 counter$count = 13186;
	#10 counter$count = 13187;
	#10 counter$count = 13188;
	#10 counter$count = 13189;
	#10 counter$count = 13190;
	#10 counter$count = 13191;
	#10 counter$count = 13192;
	#10 counter$count = 13193;
	#10 counter$count = 13194;
	#10 counter$count = 13195;
	#10 counter$count = 13196;
	#10 counter$count = 13197;
	#10 counter$count = 13198;
	#10 counter$count = 13199;
	#10 counter$count = 13200;
	#10 counter$count = 13201;
	#10 counter$count = 13202;
	#10 counter$count = 13203;
	#10 counter$count = 13204;
	#10 counter$count = 13205;
	#10 counter$count = 13206;
	#10 counter$count = 13207;
	#10 counter$count = 13208;
	#10 counter$count = 13209;
	#10 counter$count = 13210;
	#10 counter$count = 13211;
	#10 counter$count = 13212;
	#10 counter$count = 13213;
	#10 counter$count = 13214;
	#10 counter$count = 13215;
	#10 counter$count = 13216;
	#10 counter$count = 13217;
	#10 counter$count = 13218;
	#10 counter$count = 13219;
	#10 counter$count = 13220;
	#10 counter$count = 13221;
	#10 counter$count = 13222;
	#10 counter$count = 13223;
	#10 counter$count = 13224;
	#10 counter$count = 13225;
	#10 counter$count = 13226;
	#10 counter$count = 13227;
	#10 counter$count = 13228;
	#10 counter$count = 13229;
	#10 counter$count = 13230;
	#10 counter$count = 13231;
	#10 counter$count = 13232;
	#10 counter$count = 13233;
	#10 counter$count = 13234;
	#10 counter$count = 13235;
	#10 counter$count = 13236;
	#10 counter$count = 13237;
	#10 counter$count = 13238;
	#10 counter$count = 13239;
	#10 counter$count = 13240;
	#10 counter$count = 13241;
	#10 counter$count = 13242;
	#10 counter$count = 13243;
	#10 counter$count = 13244;
	#10 counter$count = 13245;
	#10 counter$count = 13246;
	#10 counter$count = 13247;
	#10 counter$count = 13248;
	#10 counter$count = 13249;
	#10 counter$count = 13250;
	#10 counter$count = 13251;
	#10 counter$count = 13252;
	#10 counter$count = 13253;
	#10 counter$count = 13254;
	#10 counter$count = 13255;
	#10 counter$count = 13256;
	#10 counter$count = 13257;
	#10 counter$count = 13258;
	#10 counter$count = 13259;
	#10 counter$count = 13260;
	#10 counter$count = 13261;
	#10 counter$count = 13262;
	#10 counter$count = 13263;
	#10 counter$count = 13264;
	#10 counter$count = 13265;
	#10 counter$count = 13266;
	#10 counter$count = 13267;
	#10 counter$count = 13268;
	#10 counter$count = 13269;
	#10 counter$count = 13270;
	#10 counter$count = 13271;
	#10 counter$count = 13272;
	#10 counter$count = 13273;
	#10 counter$count = 13274;
	#10 counter$count = 13275;
	#10 counter$count = 13276;
	#10 counter$count = 13277;
	#10 counter$count = 13278;
	#10 counter$count = 13279;
	#10 counter$count = 13280;
	#10 counter$count = 13281;
	#10 counter$count = 13282;
	#10 counter$count = 13283;
	#10 counter$count = 13284;
	#10 counter$count = 13285;
	#10 counter$count = 13286;
	#10 counter$count = 13287;
	#10 counter$count = 13288;
	#10 counter$count = 13289;
	#10 counter$count = 13290;
	#10 counter$count = 13291;
	#10 counter$count = 13292;
	#10 counter$count = 13293;
	#10 counter$count = 13294;
	#10 counter$count = 13295;
	#10 counter$count = 13296;
	#10 counter$count = 13297;
	#10 counter$count = 13298;
	#10 counter$count = 13299;
	#10 counter$count = 13300;
	#10 counter$count = 13301;
	#10 counter$count = 13302;
	#10 counter$count = 13303;
	#10 counter$count = 13304;
	#10 counter$count = 13305;
	#10 counter$count = 13306;
	#10 counter$count = 13307;
	#10 counter$count = 13308;
	#10 counter$count = 13309;
	#10 counter$count = 13310;
	#10 counter$count = 13311;
	#10 counter$count = 13312;
	#10 counter$count = 13313;
	#10 counter$count = 13314;
	#10 counter$count = 13315;
	#10 counter$count = 13316;
	#10 counter$count = 13317;
	#10 counter$count = 13318;
	#10 counter$count = 13319;
	#10 counter$count = 13320;
	#10 counter$count = 13321;
	#10 counter$count = 13322;
	#10 counter$count = 13323;
	#10 counter$count = 13324;
	#10 counter$count = 13325;
	#10 counter$count = 13326;
	#10 counter$count = 13327;
	#10 counter$count = 13328;
	#10 counter$count = 13329;
	#10 counter$count = 13330;
	#10 counter$count = 13331;
	#10 counter$count = 13332;
	#10 counter$count = 13333;
	#10 counter$count = 13334;
	#10 counter$count = 13335;
	#10 counter$count = 13336;
	#10 counter$count = 13337;
	#10 counter$count = 13338;
	#10 counter$count = 13339;
	#10 counter$count = 13340;
	#10 counter$count = 13341;
	#10 counter$count = 13342;
	#10 counter$count = 13343;
	#10 counter$count = 13344;
	#10 counter$count = 13345;
	#10 counter$count = 13346;
	#10 counter$count = 13347;
	#10 counter$count = 13348;
	#10 counter$count = 13349;
	#10 counter$count = 13350;
	#10 counter$count = 13351;
	#10 counter$count = 13352;
	#10 counter$count = 13353;
	#10 counter$count = 13354;
	#10 counter$count = 13355;
	#10 counter$count = 13356;
	#10 counter$count = 13357;
	#10 counter$count = 13358;
	#10 counter$count = 13359;
	#10 counter$count = 13360;
	#10 counter$count = 13361;
	#10 counter$count = 13362;
	#10 counter$count = 13363;
	#10 counter$count = 13364;
	#10 counter$count = 13365;
	#10 counter$count = 13366;
	#10 counter$count = 13367;
	#10 counter$count = 13368;
	#10 counter$count = 13369;
	#10 counter$count = 13370;
	#10 counter$count = 13371;
	#10 counter$count = 13372;
	#10 counter$count = 13373;
	#10 counter$count = 13374;
	#10 counter$count = 13375;
	#10 counter$count = 13376;
	#10 counter$count = 13377;
	#10 counter$count = 13378;
	#10 counter$count = 13379;
	#10 counter$count = 13380;
	#10 counter$count = 13381;
	#10 counter$count = 13382;
	#10 counter$count = 13383;
	#10 counter$count = 13384;
	#10 counter$count = 13385;
	#10 counter$count = 13386;
	#10 counter$count = 13387;
	#10 counter$count = 13388;
	#10 counter$count = 13389;
	#10 counter$count = 13390;
	#10 counter$count = 13391;
	#10 counter$count = 13392;
	#10 counter$count = 13393;
	#10 counter$count = 13394;
	#10 counter$count = 13395;
	#10 counter$count = 13396;
	#10 counter$count = 13397;
	#10 counter$count = 13398;
	#10 counter$count = 13399;
	#10 counter$count = 13400;
	#10 counter$count = 13401;
	#10 counter$count = 13402;
	#10 counter$count = 13403;
	#10 counter$count = 13404;
	#10 counter$count = 13405;
	#10 counter$count = 13406;
	#10 counter$count = 13407;
	#10 counter$count = 13408;
	#10 counter$count = 13409;
	#10 counter$count = 13410;
	#10 counter$count = 13411;
	#10 counter$count = 13412;
	#10 counter$count = 13413;
	#10 counter$count = 13414;
	#10 counter$count = 13415;
	#10 counter$count = 13416;
	#10 counter$count = 13417;
	#10 counter$count = 13418;
	#10 counter$count = 13419;
	#10 counter$count = 13420;
	#10 counter$count = 13421;
	#10 counter$count = 13422;
	#10 counter$count = 13423;
	#10 counter$count = 13424;
	#10 counter$count = 13425;
	#10 counter$count = 13426;
	#10 counter$count = 13427;
	#10 counter$count = 13428;
	#10 counter$count = 13429;
	#10 counter$count = 13430;
	#10 counter$count = 13431;
	#10 counter$count = 13432;
	#10 counter$count = 13433;
	#10 counter$count = 13434;
	#10 counter$count = 13435;
	#10 counter$count = 13436;
	#10 counter$count = 13437;
	#10 counter$count = 13438;
	#10 counter$count = 13439;
	#10 counter$count = 13440;
	#10 counter$count = 13441;
	#10 counter$count = 13442;
	#10 counter$count = 13443;
	#10 counter$count = 13444;
	#10 counter$count = 13445;
	#10 counter$count = 13446;
	#10 counter$count = 13447;
	#10 counter$count = 13448;
	#10 counter$count = 13449;
	#10 counter$count = 13450;
	#10 counter$count = 13451;
	#10 counter$count = 13452;
	#10 counter$count = 13453;
	#10 counter$count = 13454;
	#10 counter$count = 13455;
	#10 counter$count = 13456;
	#10 counter$count = 13457;
	#10 counter$count = 13458;
	#10 counter$count = 13459;
	#10 counter$count = 13460;
	#10 counter$count = 13461;
	#10 counter$count = 13462;
	#10 counter$count = 13463;
	#10 counter$count = 13464;
	#10 counter$count = 13465;
	#10 counter$count = 13466;
	#10 counter$count = 13467;
	#10 counter$count = 13468;
	#10 counter$count = 13469;
	#10 counter$count = 13470;
	#10 counter$count = 13471;
	#10 counter$count = 13472;
	#10 counter$count = 13473;
	#10 counter$count = 13474;
	#10 counter$count = 13475;
	#10 counter$count = 13476;
	#10 counter$count = 13477;
	#10 counter$count = 13478;
	#10 counter$count = 13479;
	#10 counter$count = 13480;
	#10 counter$count = 13481;
	#10 counter$count = 13482;
	#10 counter$count = 13483;
	#10 counter$count = 13484;
	#10 counter$count = 13485;
	#10 counter$count = 13486;
	#10 counter$count = 13487;
	#10 counter$count = 13488;
	#10 counter$count = 13489;
	#10 counter$count = 13490;
	#10 counter$count = 13491;
	#10 counter$count = 13492;
	#10 counter$count = 13493;
	#10 counter$count = 13494;
	#10 counter$count = 13495;
	#10 counter$count = 13496;
	#10 counter$count = 13497;
	#10 counter$count = 13498;
	#10 counter$count = 13499;
	#10 counter$count = 13500;
	#10 counter$count = 13501;
	#10 counter$count = 13502;
	#10 counter$count = 13503;
	#10 counter$count = 13504;
	#10 counter$count = 13505;
	#10 counter$count = 13506;
	#10 counter$count = 13507;
	#10 counter$count = 13508;
	#10 counter$count = 13509;
	#10 counter$count = 13510;
	#10 counter$count = 13511;
	#10 counter$count = 13512;
	#10 counter$count = 13513;
	#10 counter$count = 13514;
	#10 counter$count = 13515;
	#10 counter$count = 13516;
	#10 counter$count = 13517;
	#10 counter$count = 13518;
	#10 counter$count = 13519;
	#10 counter$count = 13520;
	#10 counter$count = 13521;
	#10 counter$count = 13522;
	#10 counter$count = 13523;
	#10 counter$count = 13524;
	#10 counter$count = 13525;
	#10 counter$count = 13526;
	#10 counter$count = 13527;
	#10 counter$count = 13528;
	#10 counter$count = 13529;
	#10 counter$count = 13530;
	#10 counter$count = 13531;
	#10 counter$count = 13532;
	#10 counter$count = 13533;
	#10 counter$count = 13534;
	#10 counter$count = 13535;
	#10 counter$count = 13536;
	#10 counter$count = 13537;
	#10 counter$count = 13538;
	#10 counter$count = 13539;
	#10 counter$count = 13540;
	#10 counter$count = 13541;
	#10 counter$count = 13542;
	#10 counter$count = 13543;
	#10 counter$count = 13544;
	#10 counter$count = 13545;
	#10 counter$count = 13546;
	#10 counter$count = 13547;
	#10 counter$count = 13548;
	#10 counter$count = 13549;
	#10 counter$count = 13550;
	#10 counter$count = 13551;
	#10 counter$count = 13552;
	#10 counter$count = 13553;
	#10 counter$count = 13554;
	#10 counter$count = 13555;
	#10 counter$count = 13556;
	#10 counter$count = 13557;
	#10 counter$count = 13558;
	#10 counter$count = 13559;
	#10 counter$count = 13560;
	#10 counter$count = 13561;
	#10 counter$count = 13562;
	#10 counter$count = 13563;
	#10 counter$count = 13564;
	#10 counter$count = 13565;
	#10 counter$count = 13566;
	#10 counter$count = 13567;
	#10 counter$count = 13568;
	#10 counter$count = 13569;
	#10 counter$count = 13570;
	#10 counter$count = 13571;
	#10 counter$count = 13572;
	#10 counter$count = 13573;
	#10 counter$count = 13574;
	#10 counter$count = 13575;
	#10 counter$count = 13576;
	#10 counter$count = 13577;
	#10 counter$count = 13578;
	#10 counter$count = 13579;
	#10 counter$count = 13580;
	#10 counter$count = 13581;
	#10 counter$count = 13582;
	#10 counter$count = 13583;
	#10 counter$count = 13584;
	#10 counter$count = 13585;
	#10 counter$count = 13586;
	#10 counter$count = 13587;
	#10 counter$count = 13588;
	#10 counter$count = 13589;
	#10 counter$count = 13590;
	#10 counter$count = 13591;
	#10 counter$count = 13592;
	#10 counter$count = 13593;
	#10 counter$count = 13594;
	#10 counter$count = 13595;
	#10 counter$count = 13596;
	#10 counter$count = 13597;
	#10 counter$count = 13598;
	#10 counter$count = 13599;
	#10 counter$count = 13600;
	#10 counter$count = 13601;
	#10 counter$count = 13602;
	#10 counter$count = 13603;
	#10 counter$count = 13604;
	#10 counter$count = 13605;
	#10 counter$count = 13606;
	#10 counter$count = 13607;
	#10 counter$count = 13608;
	#10 counter$count = 13609;
	#10 counter$count = 13610;
	#10 counter$count = 13611;
	#10 counter$count = 13612;
	#10 counter$count = 13613;
	#10 counter$count = 13614;
	#10 counter$count = 13615;
	#10 counter$count = 13616;
	#10 counter$count = 13617;
	#10 counter$count = 13618;
	#10 counter$count = 13619;
	#10 counter$count = 13620;
	#10 counter$count = 13621;
	#10 counter$count = 13622;
	#10 counter$count = 13623;
	#10 counter$count = 13624;
	#10 counter$count = 13625;
	#10 counter$count = 13626;
	#10 counter$count = 13627;
	#10 counter$count = 13628;
	#10 counter$count = 13629;
	#10 counter$count = 13630;
	#10 counter$count = 13631;
	#10 counter$count = 13632;
	#10 counter$count = 13633;
	#10 counter$count = 13634;
	#10 counter$count = 13635;
	#10 counter$count = 13636;
	#10 counter$count = 13637;
	#10 counter$count = 13638;
	#10 counter$count = 13639;
	#10 counter$count = 13640;
	#10 counter$count = 13641;
	#10 counter$count = 13642;
	#10 counter$count = 13643;
	#10 counter$count = 13644;
	#10 counter$count = 13645;
	#10 counter$count = 13646;
	#10 counter$count = 13647;
	#10 counter$count = 13648;
	#10 counter$count = 13649;
	#10 counter$count = 13650;
	#10 counter$count = 13651;
	#10 counter$count = 13652;
	#10 counter$count = 13653;
	#10 counter$count = 13654;
	#10 counter$count = 13655;
	#10 counter$count = 13656;
	#10 counter$count = 13657;
	#10 counter$count = 13658;
	#10 counter$count = 13659;
	#10 counter$count = 13660;
	#10 counter$count = 13661;
	#10 counter$count = 13662;
	#10 counter$count = 13663;
	#10 counter$count = 13664;
	#10 counter$count = 13665;
	#10 counter$count = 13666;
	#10 counter$count = 13667;
	#10 counter$count = 13668;
	#10 counter$count = 13669;
	#10 counter$count = 13670;
	#10 counter$count = 13671;
	#10 counter$count = 13672;
	#10 counter$count = 13673;
	#10 counter$count = 13674;
	#10 counter$count = 13675;
	#10 counter$count = 13676;
	#10 counter$count = 13677;
	#10 counter$count = 13678;
	#10 counter$count = 13679;
	#10 counter$count = 13680;
	#10 counter$count = 13681;
	#10 counter$count = 13682;
	#10 counter$count = 13683;
	#10 counter$count = 13684;
	#10 counter$count = 13685;
	#10 counter$count = 13686;
	#10 counter$count = 13687;
	#10 counter$count = 13688;
	#10 counter$count = 13689;
	#10 counter$count = 13690;
	#10 counter$count = 13691;
	#10 counter$count = 13692;
	#10 counter$count = 13693;
	#10 counter$count = 13694;
	#10 counter$count = 13695;
	#10 counter$count = 13696;
	#10 counter$count = 13697;
	#10 counter$count = 13698;
	#10 counter$count = 13699;
	#10 counter$count = 13700;
	#10 counter$count = 13701;
	#10 counter$count = 13702;
	#10 counter$count = 13703;
	#10 counter$count = 13704;
	#10 counter$count = 13705;
	#10 counter$count = 13706;
	#10 counter$count = 13707;
	#10 counter$count = 13708;
	#10 counter$count = 13709;
	#10 counter$count = 13710;
	#10 counter$count = 13711;
	#10 counter$count = 13712;
	#10 counter$count = 13713;
	#10 counter$count = 13714;
	#10 counter$count = 13715;
	#10 counter$count = 13716;
	#10 counter$count = 13717;
	#10 counter$count = 13718;
	#10 counter$count = 13719;
	#10 counter$count = 13720;
	#10 counter$count = 13721;
	#10 counter$count = 13722;
	#10 counter$count = 13723;
	#10 counter$count = 13724;
	#10 counter$count = 13725;
	#10 counter$count = 13726;
	#10 counter$count = 13727;
	#10 counter$count = 13728;
	#10 counter$count = 13729;
	#10 counter$count = 13730;
	#10 counter$count = 13731;
	#10 counter$count = 13732;
	#10 counter$count = 13733;
	#10 counter$count = 13734;
	#10 counter$count = 13735;
	#10 counter$count = 13736;
	#10 counter$count = 13737;
	#10 counter$count = 13738;
	#10 counter$count = 13739;
	#10 counter$count = 13740;
	#10 counter$count = 13741;
	#10 counter$count = 13742;
	#10 counter$count = 13743;
	#10 counter$count = 13744;
	#10 counter$count = 13745;
	#10 counter$count = 13746;
	#10 counter$count = 13747;
	#10 counter$count = 13748;
	#10 counter$count = 13749;
	#10 counter$count = 13750;
	#10 counter$count = 13751;
	#10 counter$count = 13752;
	#10 counter$count = 13753;
	#10 counter$count = 13754;
	#10 counter$count = 13755;
	#10 counter$count = 13756;
	#10 counter$count = 13757;
	#10 counter$count = 13758;
	#10 counter$count = 13759;
	#10 counter$count = 13760;
	#10 counter$count = 13761;
	#10 counter$count = 13762;
	#10 counter$count = 13763;
	#10 counter$count = 13764;
	#10 counter$count = 13765;
	#10 counter$count = 13766;
	#10 counter$count = 13767;
	#10 counter$count = 13768;
	#10 counter$count = 13769;
	#10 counter$count = 13770;
	#10 counter$count = 13771;
	#10 counter$count = 13772;
	#10 counter$count = 13773;
	#10 counter$count = 13774;
	#10 counter$count = 13775;
	#10 counter$count = 13776;
	#10 counter$count = 13777;
	#10 counter$count = 13778;
	#10 counter$count = 13779;
	#10 counter$count = 13780;
	#10 counter$count = 13781;
	#10 counter$count = 13782;
	#10 counter$count = 13783;
	#10 counter$count = 13784;
	#10 counter$count = 13785;
	#10 counter$count = 13786;
	#10 counter$count = 13787;
	#10 counter$count = 13788;
	#10 counter$count = 13789;
	#10 counter$count = 13790;
	#10 counter$count = 13791;
	#10 counter$count = 13792;
	#10 counter$count = 13793;
	#10 counter$count = 13794;
	#10 counter$count = 13795;
	#10 counter$count = 13796;
	#10 counter$count = 13797;
	#10 counter$count = 13798;
	#10 counter$count = 13799;
	#10 counter$count = 13800;
	#10 counter$count = 13801;
	#10 counter$count = 13802;
	#10 counter$count = 13803;
	#10 counter$count = 13804;
	#10 counter$count = 13805;
	#10 counter$count = 13806;
	#10 counter$count = 13807;
	#10 counter$count = 13808;
	#10 counter$count = 13809;
	#10 counter$count = 13810;
	#10 counter$count = 13811;
	#10 counter$count = 13812;
	#10 counter$count = 13813;
	#10 counter$count = 13814;
	#10 counter$count = 13815;
	#10 counter$count = 13816;
	#10 counter$count = 13817;
	#10 counter$count = 13818;
	#10 counter$count = 13819;
	#10 counter$count = 13820;
	#10 counter$count = 13821;
	#10 counter$count = 13822;
	#10 counter$count = 13823;
	#10 counter$count = 13824;
	#10 counter$count = 13825;
	#10 counter$count = 13826;
	#10 counter$count = 13827;
	#10 counter$count = 13828;
	#10 counter$count = 13829;
	#10 counter$count = 13830;
	#10 counter$count = 13831;
	#10 counter$count = 13832;
	#10 counter$count = 13833;
	#10 counter$count = 13834;
	#10 counter$count = 13835;
	#10 counter$count = 13836;
	#10 counter$count = 13837;
	#10 counter$count = 13838;
	#10 counter$count = 13839;
	#10 counter$count = 13840;
	#10 counter$count = 13841;
	#10 counter$count = 13842;
	#10 counter$count = 13843;
	#10 counter$count = 13844;
	#10 counter$count = 13845;
	#10 counter$count = 13846;
	#10 counter$count = 13847;
	#10 counter$count = 13848;
	#10 counter$count = 13849;
	#10 counter$count = 13850;
	#10 counter$count = 13851;
	#10 counter$count = 13852;
	#10 counter$count = 13853;
	#10 counter$count = 13854;
	#10 counter$count = 13855;
	#10 counter$count = 13856;
	#10 counter$count = 13857;
	#10 counter$count = 13858;
	#10 counter$count = 13859;
	#10 counter$count = 13860;
	#10 counter$count = 13861;
	#10 counter$count = 13862;
	#10 counter$count = 13863;
	#10 counter$count = 13864;
	#10 counter$count = 13865;
	#10 counter$count = 13866;
	#10 counter$count = 13867;
	#10 counter$count = 13868;
	#10 counter$count = 13869;
	#10 counter$count = 13870;
	#10 counter$count = 13871;
	#10 counter$count = 13872;
	#10 counter$count = 13873;
	#10 counter$count = 13874;
	#10 counter$count = 13875;
	#10 counter$count = 13876;
	#10 counter$count = 13877;
	#10 counter$count = 13878;
	#10 counter$count = 13879;
	#10 counter$count = 13880;
	#10 counter$count = 13881;
	#10 counter$count = 13882;
	#10 counter$count = 13883;
	#10 counter$count = 13884;
	#10 counter$count = 13885;
	#10 counter$count = 13886;
	#10 counter$count = 13887;
	#10 counter$count = 13888;
	#10 counter$count = 13889;
	#10 counter$count = 13890;
	#10 counter$count = 13891;
	#10 counter$count = 13892;
	#10 counter$count = 13893;
	#10 counter$count = 13894;
	#10 counter$count = 13895;
	#10 counter$count = 13896;
	#10 counter$count = 13897;
	#10 counter$count = 13898;
	#10 counter$count = 13899;
	#10 counter$count = 13900;
	#10 counter$count = 13901;
	#10 counter$count = 13902;
	#10 counter$count = 13903;
	#10 counter$count = 13904;
	#10 counter$count = 13905;
	#10 counter$count = 13906;
	#10 counter$count = 13907;
	#10 counter$count = 13908;
	#10 counter$count = 13909;
	#10 counter$count = 13910;
	#10 counter$count = 13911;
	#10 counter$count = 13912;
	#10 counter$count = 13913;
	#10 counter$count = 13914;
	#10 counter$count = 13915;
	#10 counter$count = 13916;
	#10 counter$count = 13917;
	#10 counter$count = 13918;
	#10 counter$count = 13919;
	#10 counter$count = 13920;
	#10 counter$count = 13921;
	#10 counter$count = 13922;
	#10 counter$count = 13923;
	#10 counter$count = 13924;
	#10 counter$count = 13925;
	#10 counter$count = 13926;
	#10 counter$count = 13927;
	#10 counter$count = 13928;
	#10 counter$count = 13929;
	#10 counter$count = 13930;
	#10 counter$count = 13931;
	#10 counter$count = 13932;
	#10 counter$count = 13933;
	#10 counter$count = 13934;
	#10 counter$count = 13935;
	#10 counter$count = 13936;
	#10 counter$count = 13937;
	#10 counter$count = 13938;
	#10 counter$count = 13939;
	#10 counter$count = 13940;
	#10 counter$count = 13941;
	#10 counter$count = 13942;
	#10 counter$count = 13943;
	#10 counter$count = 13944;
	#10 counter$count = 13945;
	#10 counter$count = 13946;
	#10 counter$count = 13947;
	#10 counter$count = 13948;
	#10 counter$count = 13949;
	#10 counter$count = 13950;
	#10 counter$count = 13951;
	#10 counter$count = 13952;
	#10 counter$count = 13953;
	#10 counter$count = 13954;
	#10 counter$count = 13955;
	#10 counter$count = 13956;
	#10 counter$count = 13957;
	#10 counter$count = 13958;
	#10 counter$count = 13959;
	#10 counter$count = 13960;
	#10 counter$count = 13961;
	#10 counter$count = 13962;
	#10 counter$count = 13963;
	#10 counter$count = 13964;
	#10 counter$count = 13965;
	#10 counter$count = 13966;
	#10 counter$count = 13967;
	#10 counter$count = 13968;
	#10 counter$count = 13969;
	#10 counter$count = 13970;
	#10 counter$count = 13971;
	#10 counter$count = 13972;
	#10 counter$count = 13973;
	#10 counter$count = 13974;
	#10 counter$count = 13975;
	#10 counter$count = 13976;
	#10 counter$count = 13977;
	#10 counter$count = 13978;
	#10 counter$count = 13979;
	#10 counter$count = 13980;
	#10 counter$count = 13981;
	#10 counter$count = 13982;
	#10 counter$count = 13983;
	#10 counter$count = 13984;
	#10 counter$count = 13985;
	#10 counter$count = 13986;
	#10 counter$count = 13987;
	#10 counter$count = 13988;
	#10 counter$count = 13989;
	#10 counter$count = 13990;
	#10 counter$count = 13991;
	#10 counter$count = 13992;
	#10 counter$count = 13993;
	#10 counter$count = 13994;
	#10 counter$count = 13995;
	#10 counter$count = 13996;
	#10 counter$count = 13997;
	#10 counter$count = 13998;
	#10 counter$count = 13999;
	#10 counter$count = 14000;
	#10 counter$count = 14001;
	#10 counter$count = 14002;
	#10 counter$count = 14003;
	#10 counter$count = 14004;
	#10 counter$count = 14005;
	#10 counter$count = 14006;
	#10 counter$count = 14007;
	#10 counter$count = 14008;
	#10 counter$count = 14009;
	#10 counter$count = 14010;
	#10 counter$count = 14011;
	#10 counter$count = 14012;
	#10 counter$count = 14013;
	#10 counter$count = 14014;
	#10 counter$count = 14015;
	#10 counter$count = 14016;
	#10 counter$count = 14017;
	#10 counter$count = 14018;
	#10 counter$count = 14019;
	#10 counter$count = 14020;
	#10 counter$count = 14021;
	#10 counter$count = 14022;
	#10 counter$count = 14023;
	#10 counter$count = 14024;
	#10 counter$count = 14025;
	#10 counter$count = 14026;
	#10 counter$count = 14027;
	#10 counter$count = 14028;
	#10 counter$count = 14029;
	#10 counter$count = 14030;
	#10 counter$count = 14031;
	#10 counter$count = 14032;
	#10 counter$count = 14033;
	#10 counter$count = 14034;
	#10 counter$count = 14035;
	#10 counter$count = 14036;
	#10 counter$count = 14037;
	#10 counter$count = 14038;
	#10 counter$count = 14039;
	#10 counter$count = 14040;
	#10 counter$count = 14041;
	#10 counter$count = 14042;
	#10 counter$count = 14043;
	#10 counter$count = 14044;
	#10 counter$count = 14045;
	#10 counter$count = 14046;
	#10 counter$count = 14047;
	#10 counter$count = 14048;
	#10 counter$count = 14049;
	#10 counter$count = 14050;
	#10 counter$count = 14051;
	#10 counter$count = 14052;
	#10 counter$count = 14053;
	#10 counter$count = 14054;
	#10 counter$count = 14055;
	#10 counter$count = 14056;
	#10 counter$count = 14057;
	#10 counter$count = 14058;
	#10 counter$count = 14059;
	#10 counter$count = 14060;
	#10 counter$count = 14061;
	#10 counter$count = 14062;
	#10 counter$count = 14063;
	#10 counter$count = 14064;
	#10 counter$count = 14065;
	#10 counter$count = 14066;
	#10 counter$count = 14067;
	#10 counter$count = 14068;
	#10 counter$count = 14069;
	#10 counter$count = 14070;
	#10 counter$count = 14071;
	#10 counter$count = 14072;
	#10 counter$count = 14073;
	#10 counter$count = 14074;
	#10 counter$count = 14075;
	#10 counter$count = 14076;
	#10 counter$count = 14077;
	#10 counter$count = 14078;
	#10 counter$count = 14079;
	#10 counter$count = 14080;
	#10 counter$count = 14081;
	#10 counter$count = 14082;
	#10 counter$count = 14083;
	#10 counter$count = 14084;
	#10 counter$count = 14085;
	#10 counter$count = 14086;
	#10 counter$count = 14087;
	#10 counter$count = 14088;
	#10 counter$count = 14089;
	#10 counter$count = 14090;
	#10 counter$count = 14091;
	#10 counter$count = 14092;
	#10 counter$count = 14093;
	#10 counter$count = 14094;
	#10 counter$count = 14095;
	#10 counter$count = 14096;
	#10 counter$count = 14097;
	#10 counter$count = 14098;
	#10 counter$count = 14099;
	#10 counter$count = 14100;
	#10 counter$count = 14101;
	#10 counter$count = 14102;
	#10 counter$count = 14103;
	#10 counter$count = 14104;
	#10 counter$count = 14105;
	#10 counter$count = 14106;
	#10 counter$count = 14107;
	#10 counter$count = 14108;
	#10 counter$count = 14109;
	#10 counter$count = 14110;
	#10 counter$count = 14111;
	#10 counter$count = 14112;
	#10 counter$count = 14113;
	#10 counter$count = 14114;
	#10 counter$count = 14115;
	#10 counter$count = 14116;
	#10 counter$count = 14117;
	#10 counter$count = 14118;
	#10 counter$count = 14119;
	#10 counter$count = 14120;
	#10 counter$count = 14121;
	#10 counter$count = 14122;
	#10 counter$count = 14123;
	#10 counter$count = 14124;
	#10 counter$count = 14125;
	#10 counter$count = 14126;
	#10 counter$count = 14127;
	#10 counter$count = 14128;
	#10 counter$count = 14129;
	#10 counter$count = 14130;
	#10 counter$count = 14131;
	#10 counter$count = 14132;
	#10 counter$count = 14133;
	#10 counter$count = 14134;
	#10 counter$count = 14135;
	#10 counter$count = 14136;
	#10 counter$count = 14137;
	#10 counter$count = 14138;
	#10 counter$count = 14139;
	#10 counter$count = 14140;
	#10 counter$count = 14141;
	#10 counter$count = 14142;
	#10 counter$count = 14143;
	#10 counter$count = 14144;
	#10 counter$count = 14145;
	#10 counter$count = 14146;
	#10 counter$count = 14147;
	#10 counter$count = 14148;
	#10 counter$count = 14149;
	#10 counter$count = 14150;
	#10 counter$count = 14151;
	#10 counter$count = 14152;
	#10 counter$count = 14153;
	#10 counter$count = 14154;
	#10 counter$count = 14155;
	#10 counter$count = 14156;
	#10 counter$count = 14157;
	#10 counter$count = 14158;
	#10 counter$count = 14159;
	#10 counter$count = 14160;
	#10 counter$count = 14161;
	#10 counter$count = 14162;
	#10 counter$count = 14163;
	#10 counter$count = 14164;
	#10 counter$count = 14165;
	#10 counter$count = 14166;
	#10 counter$count = 14167;
	#10 counter$count = 14168;
	#10 counter$count = 14169;
	#10 counter$count = 14170;
	#10 counter$count = 14171;
	#10 counter$count = 14172;
	#10 counter$count = 14173;
	#10 counter$count = 14174;
	#10 counter$count = 14175;
	#10 counter$count = 14176;
	#10 counter$count = 14177;
	#10 counter$count = 14178;
	#10 counter$count = 14179;
	#10 counter$count = 14180;
	#10 counter$count = 14181;
	#10 counter$count = 14182;
	#10 counter$count = 14183;
	#10 counter$count = 14184;
	#10 counter$count = 14185;
	#10 counter$count = 14186;
	#10 counter$count = 14187;
	#10 counter$count = 14188;
	#10 counter$count = 14189;
	#10 counter$count = 14190;
	#10 counter$count = 14191;
	#10 counter$count = 14192;
	#10 counter$count = 14193;
	#10 counter$count = 14194;
	#10 counter$count = 14195;
	#10 counter$count = 14196;
	#10 counter$count = 14197;
	#10 counter$count = 14198;
	#10 counter$count = 14199;
	#10 counter$count = 14200;
	#10 counter$count = 14201;
	#10 counter$count = 14202;
	#10 counter$count = 14203;
	#10 counter$count = 14204;
	#10 counter$count = 14205;
	#10 counter$count = 14206;
	#10 counter$count = 14207;
	#10 counter$count = 14208;
	#10 counter$count = 14209;
	#10 counter$count = 14210;
	#10 counter$count = 14211;
	#10 counter$count = 14212;
	#10 counter$count = 14213;
	#10 counter$count = 14214;
	#10 counter$count = 14215;
	#10 counter$count = 14216;
	#10 counter$count = 14217;
	#10 counter$count = 14218;
	#10 counter$count = 14219;
	#10 counter$count = 14220;
	#10 counter$count = 14221;
	#10 counter$count = 14222;
	#10 counter$count = 14223;
	#10 counter$count = 14224;
	#10 counter$count = 14225;
	#10 counter$count = 14226;
	#10 counter$count = 14227;
	#10 counter$count = 14228;
	#10 counter$count = 14229;
	#10 counter$count = 14230;
	#10 counter$count = 14231;
	#10 counter$count = 14232;
	#10 counter$count = 14233;
	#10 counter$count = 14234;
	#10 counter$count = 14235;
	#10 counter$count = 14236;
	#10 counter$count = 14237;
	#10 counter$count = 14238;
	#10 counter$count = 14239;
	#10 counter$count = 14240;
	#10 counter$count = 14241;
	#10 counter$count = 14242;
	#10 counter$count = 14243;
	#10 counter$count = 14244;
	#10 counter$count = 14245;
	#10 counter$count = 14246;
	#10 counter$count = 14247;
	#10 counter$count = 14248;
	#10 counter$count = 14249;
	#10 counter$count = 14250;
	#10 counter$count = 14251;
	#10 counter$count = 14252;
	#10 counter$count = 14253;
	#10 counter$count = 14254;
	#10 counter$count = 14255;
	#10 counter$count = 14256;
	#10 counter$count = 14257;
	#10 counter$count = 14258;
	#10 counter$count = 14259;
	#10 counter$count = 14260;
	#10 counter$count = 14261;
	#10 counter$count = 14262;
	#10 counter$count = 14263;
	#10 counter$count = 14264;
	#10 counter$count = 14265;
	#10 counter$count = 14266;
	#10 counter$count = 14267;
	#10 counter$count = 14268;
	#10 counter$count = 14269;
	#10 counter$count = 14270;
	#10 counter$count = 14271;
	#10 counter$count = 14272;
	#10 counter$count = 14273;
	#10 counter$count = 14274;
	#10 counter$count = 14275;
	#10 counter$count = 14276;
	#10 counter$count = 14277;
	#10 counter$count = 14278;
	#10 counter$count = 14279;
	#10 counter$count = 14280;
	#10 counter$count = 14281;
	#10 counter$count = 14282;
	#10 counter$count = 14283;
	#10 counter$count = 14284;
	#10 counter$count = 14285;
	#10 counter$count = 14286;
	#10 counter$count = 14287;
	#10 counter$count = 14288;
	#10 counter$count = 14289;
	#10 counter$count = 14290;
	#10 counter$count = 14291;
	#10 counter$count = 14292;
	#10 counter$count = 14293;
	#10 counter$count = 14294;
	#10 counter$count = 14295;
	#10 counter$count = 14296;
	#10 counter$count = 14297;
	#10 counter$count = 14298;
	#10 counter$count = 14299;
	#10 counter$count = 14300;
	#10 counter$count = 14301;
	#10 counter$count = 14302;
	#10 counter$count = 14303;
	#10 counter$count = 14304;
	#10 counter$count = 14305;
	#10 counter$count = 14306;
	#10 counter$count = 14307;
	#10 counter$count = 14308;
	#10 counter$count = 14309;
	#10 counter$count = 14310;
	#10 counter$count = 14311;
	#10 counter$count = 14312;
	#10 counter$count = 14313;
	#10 counter$count = 14314;
	#10 counter$count = 14315;
	#10 counter$count = 14316;
	#10 counter$count = 14317;
	#10 counter$count = 14318;
	#10 counter$count = 14319;
	#10 counter$count = 14320;
	#10 counter$count = 14321;
	#10 counter$count = 14322;
	#10 counter$count = 14323;
	#10 counter$count = 14324;
	#10 counter$count = 14325;
	#10 counter$count = 14326;
	#10 counter$count = 14327;
	#10 counter$count = 14328;
	#10 counter$count = 14329;
	#10 counter$count = 14330;
	#10 counter$count = 14331;
	#10 counter$count = 14332;
	#10 counter$count = 14333;
	#10 counter$count = 14334;
	#10 counter$count = 14335;
	#10 counter$count = 14336;
	#10 counter$count = 14337;
	#10 counter$count = 14338;
	#10 counter$count = 14339;
	#10 counter$count = 14340;
	#10 counter$count = 14341;
	#10 counter$count = 14342;
	#10 counter$count = 14343;
	#10 counter$count = 14344;
	#10 counter$count = 14345;
	#10 counter$count = 14346;
	#10 counter$count = 14347;
	#10 counter$count = 14348;
	#10 counter$count = 14349;
	#10 counter$count = 14350;
	#10 counter$count = 14351;
	#10 counter$count = 14352;
	#10 counter$count = 14353;
	#10 counter$count = 14354;
	#10 counter$count = 14355;
	#10 counter$count = 14356;
	#10 counter$count = 14357;
	#10 counter$count = 14358;
	#10 counter$count = 14359;
	#10 counter$count = 14360;
	#10 counter$count = 14361;
	#10 counter$count = 14362;
	#10 counter$count = 14363;
	#10 counter$count = 14364;
	#10 counter$count = 14365;
	#10 counter$count = 14366;
	#10 counter$count = 14367;
	#10 counter$count = 14368;
	#10 counter$count = 14369;
	#10 counter$count = 14370;
	#10 counter$count = 14371;
	#10 counter$count = 14372;
	#10 counter$count = 14373;
	#10 counter$count = 14374;
	#10 counter$count = 14375;
	#10 counter$count = 14376;
	#10 counter$count = 14377;
	#10 counter$count = 14378;
	#10 counter$count = 14379;
	#10 counter$count = 14380;
	#10 counter$count = 14381;
	#10 counter$count = 14382;
	#10 counter$count = 14383;
	#10 counter$count = 14384;
	#10 counter$count = 14385;
	#10 counter$count = 14386;
	#10 counter$count = 14387;
	#10 counter$count = 14388;
	#10 counter$count = 14389;
	#10 counter$count = 14390;
	#10 counter$count = 14391;
	#10 counter$count = 14392;
	#10 counter$count = 14393;
	#10 counter$count = 14394;
	#10 counter$count = 14395;
	#10 counter$count = 14396;
	#10 counter$count = 14397;
	#10 counter$count = 14398;
	#10 counter$count = 14399;
	#10 counter$count = 14400;
	#10 counter$count = 14401;
	#10 counter$count = 14402;
	#10 counter$count = 14403;
	#10 counter$count = 14404;
	#10 counter$count = 14405;
	#10 counter$count = 14406;
	#10 counter$count = 14407;
	#10 counter$count = 14408;
	#10 counter$count = 14409;
	#10 counter$count = 14410;
	#10 counter$count = 14411;
	#10 counter$count = 14412;
	#10 counter$count = 14413;
	#10 counter$count = 14414;
	#10 counter$count = 14415;
	#10 counter$count = 14416;
	#10 counter$count = 14417;
	#10 counter$count = 14418;
	#10 counter$count = 14419;
	#10 counter$count = 14420;
	#10 counter$count = 14421;
	#10 counter$count = 14422;
	#10 counter$count = 14423;
	#10 counter$count = 14424;
	#10 counter$count = 14425;
	#10 counter$count = 14426;
	#10 counter$count = 14427;
	#10 counter$count = 14428;
	#10 counter$count = 14429;
	#10 counter$count = 14430;
	#10 counter$count = 14431;
	#10 counter$count = 14432;
	#10 counter$count = 14433;
	#10 counter$count = 14434;
	#10 counter$count = 14435;
	#10 counter$count = 14436;
	#10 counter$count = 14437;
	#10 counter$count = 14438;
	#10 counter$count = 14439;
	#10 counter$count = 14440;
	#10 counter$count = 14441;
	#10 counter$count = 14442;
	#10 counter$count = 14443;
	#10 counter$count = 14444;
	#10 counter$count = 14445;
	#10 counter$count = 14446;
	#10 counter$count = 14447;
	#10 counter$count = 14448;
	#10 counter$count = 14449;
	#10 counter$count = 14450;
	#10 counter$count = 14451;
	#10 counter$count = 14452;
	#10 counter$count = 14453;
	#10 counter$count = 14454;
	#10 counter$count = 14455;
	#10 counter$count = 14456;
	#10 counter$count = 14457;
	#10 counter$count = 14458;
	#10 counter$count = 14459;
	#10 counter$count = 14460;
	#10 counter$count = 14461;
	#10 counter$count = 14462;
	#10 counter$count = 14463;
	#10 counter$count = 14464;
	#10 counter$count = 14465;
	#10 counter$count = 14466;
	#10 counter$count = 14467;
	#10 counter$count = 14468;
	#10 counter$count = 14469;
	#10 counter$count = 14470;
	#10 counter$count = 14471;
	#10 counter$count = 14472;
	#10 counter$count = 14473;
	#10 counter$count = 14474;
	#10 counter$count = 14475;
	#10 counter$count = 14476;
	#10 counter$count = 14477;
	#10 counter$count = 14478;
	#10 counter$count = 14479;
	#10 counter$count = 14480;
	#10 counter$count = 14481;
	#10 counter$count = 14482;
	#10 counter$count = 14483;
	#10 counter$count = 14484;
	#10 counter$count = 14485;
	#10 counter$count = 14486;
	#10 counter$count = 14487;
	#10 counter$count = 14488;
	#10 counter$count = 14489;
	#10 counter$count = 14490;
	#10 counter$count = 14491;
	#10 counter$count = 14492;
	#10 counter$count = 14493;
	#10 counter$count = 14494;
	#10 counter$count = 14495;
	#10 counter$count = 14496;
	#10 counter$count = 14497;
	#10 counter$count = 14498;
	#10 counter$count = 14499;
	#10 counter$count = 14500;
	#10 counter$count = 14501;
	#10 counter$count = 14502;
	#10 counter$count = 14503;
	#10 counter$count = 14504;
	#10 counter$count = 14505;
	#10 counter$count = 14506;
	#10 counter$count = 14507;
	#10 counter$count = 14508;
	#10 counter$count = 14509;
	#10 counter$count = 14510;
	#10 counter$count = 14511;
	#10 counter$count = 14512;
	#10 counter$count = 14513;
	#10 counter$count = 14514;
	#10 counter$count = 14515;
	#10 counter$count = 14516;
	#10 counter$count = 14517;
	#10 counter$count = 14518;
	#10 counter$count = 14519;
	#10 counter$count = 14520;
	#10 counter$count = 14521;
	#10 counter$count = 14522;
	#10 counter$count = 14523;
	#10 counter$count = 14524;
	#10 counter$count = 14525;
	#10 counter$count = 14526;
	#10 counter$count = 14527;
	#10 counter$count = 14528;
	#10 counter$count = 14529;
	#10 counter$count = 14530;
	#10 counter$count = 14531;
	#10 counter$count = 14532;
	#10 counter$count = 14533;
	#10 counter$count = 14534;
	#10 counter$count = 14535;
	#10 counter$count = 14536;
	#10 counter$count = 14537;
	#10 counter$count = 14538;
	#10 counter$count = 14539;
	#10 counter$count = 14540;
	#10 counter$count = 14541;
	#10 counter$count = 14542;
	#10 counter$count = 14543;
	#10 counter$count = 14544;
	#10 counter$count = 14545;
	#10 counter$count = 14546;
	#10 counter$count = 14547;
	#10 counter$count = 14548;
	#10 counter$count = 14549;
	#10 counter$count = 14550;
	#10 counter$count = 14551;
	#10 counter$count = 14552;
	#10 counter$count = 14553;
	#10 counter$count = 14554;
	#10 counter$count = 14555;
	#10 counter$count = 14556;
	#10 counter$count = 14557;
	#10 counter$count = 14558;
	#10 counter$count = 14559;
	#10 counter$count = 14560;
	#10 counter$count = 14561;
	#10 counter$count = 14562;
	#10 counter$count = 14563;
	#10 counter$count = 14564;
	#10 counter$count = 14565;
	#10 counter$count = 14566;
	#10 counter$count = 14567;
	#10 counter$count = 14568;
	#10 counter$count = 14569;
	#10 counter$count = 14570;
	#10 counter$count = 14571;
	#10 counter$count = 14572;
	#10 counter$count = 14573;
	#10 counter$count = 14574;
	#10 counter$count = 14575;
	#10 counter$count = 14576;
	#10 counter$count = 14577;
	#10 counter$count = 14578;
	#10 counter$count = 14579;
	#10 counter$count = 14580;
	#10 counter$count = 14581;
	#10 counter$count = 14582;
	#10 counter$count = 14583;
	#10 counter$count = 14584;
	#10 counter$count = 14585;
	#10 counter$count = 14586;
	#10 counter$count = 14587;
	#10 counter$count = 14588;
	#10 counter$count = 14589;
	#10 counter$count = 14590;
	#10 counter$count = 14591;
	#10 counter$count = 14592;
	#10 counter$count = 14593;
	#10 counter$count = 14594;
	#10 counter$count = 14595;
	#10 counter$count = 14596;
	#10 counter$count = 14597;
	#10 counter$count = 14598;
	#10 counter$count = 14599;
	#10 counter$count = 14600;
	#10 counter$count = 14601;
	#10 counter$count = 14602;
	#10 counter$count = 14603;
	#10 counter$count = 14604;
	#10 counter$count = 14605;
	#10 counter$count = 14606;
	#10 counter$count = 14607;
	#10 counter$count = 14608;
	#10 counter$count = 14609;
	#10 counter$count = 14610;
	#10 counter$count = 14611;
	#10 counter$count = 14612;
	#10 counter$count = 14613;
	#10 counter$count = 14614;
	#10 counter$count = 14615;
	#10 counter$count = 14616;
	#10 counter$count = 14617;
	#10 counter$count = 14618;
	#10 counter$count = 14619;
	#10 counter$count = 14620;
	#10 counter$count = 14621;
	#10 counter$count = 14622;
	#10 counter$count = 14623;
	#10 counter$count = 14624;
	#10 counter$count = 14625;
	#10 counter$count = 14626;
	#10 counter$count = 14627;
	#10 counter$count = 14628;
	#10 counter$count = 14629;
	#10 counter$count = 14630;
	#10 counter$count = 14631;
	#10 counter$count = 14632;
	#10 counter$count = 14633;
	#10 counter$count = 14634;
	#10 counter$count = 14635;
	#10 counter$count = 14636;
	#10 counter$count = 14637;
	#10 counter$count = 14638;
	#10 counter$count = 14639;
	#10 counter$count = 14640;
	#10 counter$count = 14641;
	#10 counter$count = 14642;
	#10 counter$count = 14643;
	#10 counter$count = 14644;
	#10 counter$count = 14645;
	#10 counter$count = 14646;
	#10 counter$count = 14647;
	#10 counter$count = 14648;
	#10 counter$count = 14649;
	#10 counter$count = 14650;
	#10 counter$count = 14651;
	#10 counter$count = 14652;
	#10 counter$count = 14653;
	#10 counter$count = 14654;
	#10 counter$count = 14655;
	#10 counter$count = 14656;
	#10 counter$count = 14657;
	#10 counter$count = 14658;
	#10 counter$count = 14659;
	#10 counter$count = 14660;
	#10 counter$count = 14661;
	#10 counter$count = 14662;
	#10 counter$count = 14663;
	#10 counter$count = 14664;
	#10 counter$count = 14665;
	#10 counter$count = 14666;
	#10 counter$count = 14667;
	#10 counter$count = 14668;
	#10 counter$count = 14669;
	#10 counter$count = 14670;
	#10 counter$count = 14671;
	#10 counter$count = 14672;
	#10 counter$count = 14673;
	#10 counter$count = 14674;
	#10 counter$count = 14675;
	#10 counter$count = 14676;
	#10 counter$count = 14677;
	#10 counter$count = 14678;
	#10 counter$count = 14679;
	#10 counter$count = 14680;
	#10 counter$count = 14681;
	#10 counter$count = 14682;
	#10 counter$count = 14683;
	#10 counter$count = 14684;
	#10 counter$count = 14685;
	#10 counter$count = 14686;
	#10 counter$count = 14687;
	#10 counter$count = 14688;
	#10 counter$count = 14689;
	#10 counter$count = 14690;
	#10 counter$count = 14691;
	#10 counter$count = 14692;
	#10 counter$count = 14693;
	#10 counter$count = 14694;
	#10 counter$count = 14695;
	#10 counter$count = 14696;
	#10 counter$count = 14697;
	#10 counter$count = 14698;
	#10 counter$count = 14699;
	#10 counter$count = 14700;
	#10 counter$count = 14701;
	#10 counter$count = 14702;
	#10 counter$count = 14703;
	#10 counter$count = 14704;
	#10 counter$count = 14705;
	#10 counter$count = 14706;
	#10 counter$count = 14707;
	#10 counter$count = 14708;
	#10 counter$count = 14709;
	#10 counter$count = 14710;
	#10 counter$count = 14711;
	#10 counter$count = 14712;
	#10 counter$count = 14713;
	#10 counter$count = 14714;
	#10 counter$count = 14715;
	#10 counter$count = 14716;
	#10 counter$count = 14717;
	#10 counter$count = 14718;
	#10 counter$count = 14719;
	#10 counter$count = 14720;
	#10 counter$count = 14721;
	#10 counter$count = 14722;
	#10 counter$count = 14723;
	#10 counter$count = 14724;
	#10 counter$count = 14725;
	#10 counter$count = 14726;
	#10 counter$count = 14727;
	#10 counter$count = 14728;
	#10 counter$count = 14729;
	#10 counter$count = 14730;
	#10 counter$count = 14731;
	#10 counter$count = 14732;
	#10 counter$count = 14733;
	#10 counter$count = 14734;
	#10 counter$count = 14735;
	#10 counter$count = 14736;
	#10 counter$count = 14737;
	#10 counter$count = 14738;
	#10 counter$count = 14739;
	#10 counter$count = 14740;
	#10 counter$count = 14741;
	#10 counter$count = 14742;
	#10 counter$count = 14743;
	#10 counter$count = 14744;
	#10 counter$count = 14745;
	#10 counter$count = 14746;
	#10 counter$count = 14747;
	#10 counter$count = 14748;
	#10 counter$count = 14749;
	#10 counter$count = 14750;
	#10 counter$count = 14751;
	#10 counter$count = 14752;
	#10 counter$count = 14753;
	#10 counter$count = 14754;
	#10 counter$count = 14755;
	#10 counter$count = 14756;
	#10 counter$count = 14757;
	#10 counter$count = 14758;
	#10 counter$count = 14759;
	#10 counter$count = 14760;
	#10 counter$count = 14761;
	#10 counter$count = 14762;
	#10 counter$count = 14763;
	#10 counter$count = 14764;
	#10 counter$count = 14765;
	#10 counter$count = 14766;
	#10 counter$count = 14767;
	#10 counter$count = 14768;
	#10 counter$count = 14769;
	#10 counter$count = 14770;
	#10 counter$count = 14771;
	#10 counter$count = 14772;
	#10 counter$count = 14773;
	#10 counter$count = 14774;
	#10 counter$count = 14775;
	#10 counter$count = 14776;
	#10 counter$count = 14777;
	#10 counter$count = 14778;
	#10 counter$count = 14779;
	#10 counter$count = 14780;
	#10 counter$count = 14781;
	#10 counter$count = 14782;
	#10 counter$count = 14783;
	#10 counter$count = 14784;
	#10 counter$count = 14785;
	#10 counter$count = 14786;
	#10 counter$count = 14787;
	#10 counter$count = 14788;
	#10 counter$count = 14789;
	#10 counter$count = 14790;
	#10 counter$count = 14791;
	#10 counter$count = 14792;
	#10 counter$count = 14793;
	#10 counter$count = 14794;
	#10 counter$count = 14795;
	#10 counter$count = 14796;
	#10 counter$count = 14797;
	#10 counter$count = 14798;
	#10 counter$count = 14799;
	#10 counter$count = 14800;
	#10 counter$count = 14801;
	#10 counter$count = 14802;
	#10 counter$count = 14803;
	#10 counter$count = 14804;
	#10 counter$count = 14805;
	#10 counter$count = 14806;
	#10 counter$count = 14807;
	#10 counter$count = 14808;
	#10 counter$count = 14809;
	#10 counter$count = 14810;
	#10 counter$count = 14811;
	#10 counter$count = 14812;
	#10 counter$count = 14813;
	#10 counter$count = 14814;
	#10 counter$count = 14815;
	#10 counter$count = 14816;
	#10 counter$count = 14817;
	#10 counter$count = 14818;
	#10 counter$count = 14819;
	#10 counter$count = 14820;
	#10 counter$count = 14821;
	#10 counter$count = 14822;
	#10 counter$count = 14823;
	#10 counter$count = 14824;
	#10 counter$count = 14825;
	#10 counter$count = 14826;
	#10 counter$count = 14827;
	#10 counter$count = 14828;
	#10 counter$count = 14829;
	#10 counter$count = 14830;
	#10 counter$count = 14831;
	#10 counter$count = 14832;
	#10 counter$count = 14833;
	#10 counter$count = 14834;
	#10 counter$count = 14835;
	#10 counter$count = 14836;
	#10 counter$count = 14837;
	#10 counter$count = 14838;
	#10 counter$count = 14839;
	#10 counter$count = 14840;
	#10 counter$count = 14841;
	#10 counter$count = 14842;
	#10 counter$count = 14843;
	#10 counter$count = 14844;
	#10 counter$count = 14845;
	#10 counter$count = 14846;
	#10 counter$count = 14847;
	#10 counter$count = 14848;
	#10 counter$count = 14849;
	#10 counter$count = 14850;
	#10 counter$count = 14851;
	#10 counter$count = 14852;
	#10 counter$count = 14853;
	#10 counter$count = 14854;
	#10 counter$count = 14855;
	#10 counter$count = 14856;
	#10 counter$count = 14857;
	#10 counter$count = 14858;
	#10 counter$count = 14859;
	#10 counter$count = 14860;
	#10 counter$count = 14861;
	#10 counter$count = 14862;
	#10 counter$count = 14863;
	#10 counter$count = 14864;
	#10 counter$count = 14865;
	#10 counter$count = 14866;
	#10 counter$count = 14867;
	#10 counter$count = 14868;
	#10 counter$count = 14869;
	#10 counter$count = 14870;
	#10 counter$count = 14871;
	#10 counter$count = 14872;
	#10 counter$count = 14873;
	#10 counter$count = 14874;
	#10 counter$count = 14875;
	#10 counter$count = 14876;
	#10 counter$count = 14877;
	#10 counter$count = 14878;
	#10 counter$count = 14879;
	#10 counter$count = 14880;
	#10 counter$count = 14881;
	#10 counter$count = 14882;
	#10 counter$count = 14883;
	#10 counter$count = 14884;
	#10 counter$count = 14885;
	#10 counter$count = 14886;
	#10 counter$count = 14887;
	#10 counter$count = 14888;
	#10 counter$count = 14889;
	#10 counter$count = 14890;
	#10 counter$count = 14891;
	#10 counter$count = 14892;
	#10 counter$count = 14893;
	#10 counter$count = 14894;
	#10 counter$count = 14895;
	#10 counter$count = 14896;
	#10 counter$count = 14897;
	#10 counter$count = 14898;
	#10 counter$count = 14899;
	#10 counter$count = 14900;
	#10 counter$count = 14901;
	#10 counter$count = 14902;
	#10 counter$count = 14903;
	#10 counter$count = 14904;
	#10 counter$count = 14905;
	#10 counter$count = 14906;
	#10 counter$count = 14907;
	#10 counter$count = 14908;
	#10 counter$count = 14909;
	#10 counter$count = 14910;
	#10 counter$count = 14911;
	#10 counter$count = 14912;
	#10 counter$count = 14913;
	#10 counter$count = 14914;
	#10 counter$count = 14915;
	#10 counter$count = 14916;
	#10 counter$count = 14917;
	#10 counter$count = 14918;
	#10 counter$count = 14919;
	#10 counter$count = 14920;
	#10 counter$count = 14921;
	#10 counter$count = 14922;
	#10 counter$count = 14923;
	#10 counter$count = 14924;
	#10 counter$count = 14925;
	#10 counter$count = 14926;
	#10 counter$count = 14927;
	#10 counter$count = 14928;
	#10 counter$count = 14929;
	#10 counter$count = 14930;
	#10 counter$count = 14931;
	#10 counter$count = 14932;
	#10 counter$count = 14933;
	#10 counter$count = 14934;
	#10 counter$count = 14935;
	#10 counter$count = 14936;
	#10 counter$count = 14937;
	#10 counter$count = 14938;
	#10 counter$count = 14939;
	#10 counter$count = 14940;
	#10 counter$count = 14941;
	#10 counter$count = 14942;
	#10 counter$count = 14943;
	#10 counter$count = 14944;
	#10 counter$count = 14945;
	#10 counter$count = 14946;
	#10 counter$count = 14947;
	#10 counter$count = 14948;
	#10 counter$count = 14949;
	#10 counter$count = 14950;
	#10 counter$count = 14951;
	#10 counter$count = 14952;
	#10 counter$count = 14953;
	#10 counter$count = 14954;
	#10 counter$count = 14955;
	#10 counter$count = 14956;
	#10 counter$count = 14957;
	#10 counter$count = 14958;
	#10 counter$count = 14959;
	#10 counter$count = 14960;
	#10 counter$count = 14961;
	#10 counter$count = 14962;
	#10 counter$count = 14963;
	#10 counter$count = 14964;
	#10 counter$count = 14965;
	#10 counter$count = 14966;
	#10 counter$count = 14967;
	#10 counter$count = 14968;
	#10 counter$count = 14969;
	#10 counter$count = 14970;
	#10 counter$count = 14971;
	#10 counter$count = 14972;
	#10 counter$count = 14973;
	#10 counter$count = 14974;
	#10 counter$count = 14975;
	#10 counter$count = 14976;
	#10 counter$count = 14977;
	#10 counter$count = 14978;
	#10 counter$count = 14979;
	#10 counter$count = 14980;
	#10 counter$count = 14981;
	#10 counter$count = 14982;
	#10 counter$count = 14983;
	#10 counter$count = 14984;
	#10 counter$count = 14985;
	#10 counter$count = 14986;
	#10 counter$count = 14987;
	#10 counter$count = 14988;
	#10 counter$count = 14989;
	#10 counter$count = 14990;
	#10 counter$count = 14991;
	#10 counter$count = 14992;
	#10 counter$count = 14993;
	#10 counter$count = 14994;
	#10 counter$count = 14995;
	#10 counter$count = 14996;
	#10 counter$count = 14997;
	#10 counter$count = 14998;
	#10 counter$count = 14999;
	#10 counter$count = 15000;
	#10 counter$count = 15001;
	#10 counter$count = 15002;
	#10 counter$count = 15003;
	#10 counter$count = 15004;
	#10 counter$count = 15005;
	#10 counter$count = 15006;
	#10 counter$count = 15007;
	#10 counter$count = 15008;
	#10 counter$count = 15009;
	#10 counter$count = 15010;
	#10 counter$count = 15011;
	#10 counter$count = 15012;
	#10 counter$count = 15013;
	#10 counter$count = 15014;
	#10 counter$count = 15015;
	#10 counter$count = 15016;
	#10 counter$count = 15017;
	#10 counter$count = 15018;
	#10 counter$count = 15019;
	#10 counter$count = 15020;
	#10 counter$count = 15021;
	#10 counter$count = 15022;
	#10 counter$count = 15023;
	#10 counter$count = 15024;
	#10 counter$count = 15025;
	#10 counter$count = 15026;
	#10 counter$count = 15027;
	#10 counter$count = 15028;
	#10 counter$count = 15029;
	#10 counter$count = 15030;
	#10 counter$count = 15031;
	#10 counter$count = 15032;
	#10 counter$count = 15033;
	#10 counter$count = 15034;
	#10 counter$count = 15035;
	#10 counter$count = 15036;
	#10 counter$count = 15037;
	#10 counter$count = 15038;
	#10 counter$count = 15039;
	#10 counter$count = 15040;
	#10 counter$count = 15041;
	#10 counter$count = 15042;
	#10 counter$count = 15043;
	#10 counter$count = 15044;
	#10 counter$count = 15045;
	#10 counter$count = 15046;
	#10 counter$count = 15047;
	#10 counter$count = 15048;
	#10 counter$count = 15049;
	#10 counter$count = 15050;
	#10 counter$count = 15051;
	#10 counter$count = 15052;
	#10 counter$count = 15053;
	#10 counter$count = 15054;
	#10 counter$count = 15055;
	#10 counter$count = 15056;
	#10 counter$count = 15057;
	#10 counter$count = 15058;
	#10 counter$count = 15059;
	#10 counter$count = 15060;
	#10 counter$count = 15061;
	#10 counter$count = 15062;
	#10 counter$count = 15063;
	#10 counter$count = 15064;
	#10 counter$count = 15065;
	#10 counter$count = 15066;
	#10 counter$count = 15067;
	#10 counter$count = 15068;
	#10 counter$count = 15069;
	#10 counter$count = 15070;
	#10 counter$count = 15071;
	#10 counter$count = 15072;
	#10 counter$count = 15073;
	#10 counter$count = 15074;
	#10 counter$count = 15075;
	#10 counter$count = 15076;
	#10 counter$count = 15077;
	#10 counter$count = 15078;
	#10 counter$count = 15079;
	#10 counter$count = 15080;
	#10 counter$count = 15081;
	#10 counter$count = 15082;
	#10 counter$count = 15083;
	#10 counter$count = 15084;
	#10 counter$count = 15085;
	#10 counter$count = 15086;
	#10 counter$count = 15087;
	#10 counter$count = 15088;
	#10 counter$count = 15089;
	#10 counter$count = 15090;
	#10 counter$count = 15091;
	#10 counter$count = 15092;
	#10 counter$count = 15093;
	#10 counter$count = 15094;
	#10 counter$count = 15095;
	#10 counter$count = 15096;
	#10 counter$count = 15097;
	#10 counter$count = 15098;
	#10 counter$count = 15099;
	#10 counter$count = 15100;
	#10 counter$count = 15101;
	#10 counter$count = 15102;
	#10 counter$count = 15103;
	#10 counter$count = 15104;
	#10 counter$count = 15105;
	#10 counter$count = 15106;
	#10 counter$count = 15107;
	#10 counter$count = 15108;
	#10 counter$count = 15109;
	#10 counter$count = 15110;
	#10 counter$count = 15111;
	#10 counter$count = 15112;
	#10 counter$count = 15113;
	#10 counter$count = 15114;
	#10 counter$count = 15115;
	#10 counter$count = 15116;
	#10 counter$count = 15117;
	#10 counter$count = 15118;
	#10 counter$count = 15119;
	#10 counter$count = 15120;
	#10 counter$count = 15121;
	#10 counter$count = 15122;
	#10 counter$count = 15123;
	#10 counter$count = 15124;
	#10 counter$count = 15125;
	#10 counter$count = 15126;
	#10 counter$count = 15127;
	#10 counter$count = 15128;
	#10 counter$count = 15129;
	#10 counter$count = 15130;
	#10 counter$count = 15131;
	#10 counter$count = 15132;
	#10 counter$count = 15133;
	#10 counter$count = 15134;
	#10 counter$count = 15135;
	#10 counter$count = 15136;
	#10 counter$count = 15137;
	#10 counter$count = 15138;
	#10 counter$count = 15139;
	#10 counter$count = 15140;
	#10 counter$count = 15141;
	#10 counter$count = 15142;
	#10 counter$count = 15143;
	#10 counter$count = 15144;
	#10 counter$count = 15145;
	#10 counter$count = 15146;
	#10 counter$count = 15147;
	#10 counter$count = 15148;
	#10 counter$count = 15149;
	#10 counter$count = 15150;
	#10 counter$count = 15151;
	#10 counter$count = 15152;
	#10 counter$count = 15153;
	#10 counter$count = 15154;
	#10 counter$count = 15155;
	#10 counter$count = 15156;
	#10 counter$count = 15157;
	#10 counter$count = 15158;
	#10 counter$count = 15159;
	#10 counter$count = 15160;
	#10 counter$count = 15161;
	#10 counter$count = 15162;
	#10 counter$count = 15163;
	#10 counter$count = 15164;
	#10 counter$count = 15165;
	#10 counter$count = 15166;
	#10 counter$count = 15167;
	#10 counter$count = 15168;
	#10 counter$count = 15169;
	#10 counter$count = 15170;
	#10 counter$count = 15171;
	#10 counter$count = 15172;
	#10 counter$count = 15173;
	#10 counter$count = 15174;
	#10 counter$count = 15175;
	#10 counter$count = 15176;
	#10 counter$count = 15177;
	#10 counter$count = 15178;
	#10 counter$count = 15179;
	#10 counter$count = 15180;
	#10 counter$count = 15181;
	#10 counter$count = 15182;
	#10 counter$count = 15183;
	#10 counter$count = 15184;
	#10 counter$count = 15185;
	#10 counter$count = 15186;
	#10 counter$count = 15187;
	#10 counter$count = 15188;
	#10 counter$count = 15189;
	#10 counter$count = 15190;
	#10 counter$count = 15191;
	#10 counter$count = 15192;
	#10 counter$count = 15193;
	#10 counter$count = 15194;
	#10 counter$count = 15195;
	#10 counter$count = 15196;
	#10 counter$count = 15197;
	#10 counter$count = 15198;
	#10 counter$count = 15199;
	#10 counter$count = 15200;
	#10 counter$count = 15201;
	#10 counter$count = 15202;
	#10 counter$count = 15203;
	#10 counter$count = 15204;
	#10 counter$count = 15205;
	#10 counter$count = 15206;
	#10 counter$count = 15207;
	#10 counter$count = 15208;
	#10 counter$count = 15209;
	#10 counter$count = 15210;
	#10 counter$count = 15211;
	#10 counter$count = 15212;
	#10 counter$count = 15213;
	#10 counter$count = 15214;
	#10 counter$count = 15215;
	#10 counter$count = 15216;
	#10 counter$count = 15217;
	#10 counter$count = 15218;
	#10 counter$count = 15219;
	#10 counter$count = 15220;
	#10 counter$count = 15221;
	#10 counter$count = 15222;
	#10 counter$count = 15223;
	#10 counter$count = 15224;
	#10 counter$count = 15225;
	#10 counter$count = 15226;
	#10 counter$count = 15227;
	#10 counter$count = 15228;
	#10 counter$count = 15229;
	#10 counter$count = 15230;
	#10 counter$count = 15231;
	#10 counter$count = 15232;
	#10 counter$count = 15233;
	#10 counter$count = 15234;
	#10 counter$count = 15235;
	#10 counter$count = 15236;
	#10 counter$count = 15237;
	#10 counter$count = 15238;
	#10 counter$count = 15239;
	#10 counter$count = 15240;
	#10 counter$count = 15241;
	#10 counter$count = 15242;
	#10 counter$count = 15243;
	#10 counter$count = 15244;
	#10 counter$count = 15245;
	#10 counter$count = 15246;
	#10 counter$count = 15247;
	#10 counter$count = 15248;
	#10 counter$count = 15249;
	#10 counter$count = 15250;
	#10 counter$count = 15251;
	#10 counter$count = 15252;
	#10 counter$count = 15253;
	#10 counter$count = 15254;
	#10 counter$count = 15255;
	#10 counter$count = 15256;
	#10 counter$count = 15257;
	#10 counter$count = 15258;
	#10 counter$count = 15259;
	#10 counter$count = 15260;
	#10 counter$count = 15261;
	#10 counter$count = 15262;
	#10 counter$count = 15263;
	#10 counter$count = 15264;
	#10 counter$count = 15265;
	#10 counter$count = 15266;
	#10 counter$count = 15267;
	#10 counter$count = 15268;
	#10 counter$count = 15269;
	#10 counter$count = 15270;
	#10 counter$count = 15271;
	#10 counter$count = 15272;
	#10 counter$count = 15273;
	#10 counter$count = 15274;
	#10 counter$count = 15275;
	#10 counter$count = 15276;
	#10 counter$count = 15277;
	#10 counter$count = 15278;
	#10 counter$count = 15279;
	#10 counter$count = 15280;
	#10 counter$count = 15281;
	#10 counter$count = 15282;
	#10 counter$count = 15283;
	#10 counter$count = 15284;
	#10 counter$count = 15285;
	#10 counter$count = 15286;
	#10 counter$count = 15287;
	#10 counter$count = 15288;
	#10 counter$count = 15289;
	#10 counter$count = 15290;
	#10 counter$count = 15291;
	#10 counter$count = 15292;
	#10 counter$count = 15293;
	#10 counter$count = 15294;
	#10 counter$count = 15295;
	#10 counter$count = 15296;
	#10 counter$count = 15297;
	#10 counter$count = 15298;
	#10 counter$count = 15299;
	#10 counter$count = 15300;
	#10 counter$count = 15301;
	#10 counter$count = 15302;
	#10 counter$count = 15303;
	#10 counter$count = 15304;
	#10 counter$count = 15305;
	#10 counter$count = 15306;
	#10 counter$count = 15307;
	#10 counter$count = 15308;
	#10 counter$count = 15309;
	#10 counter$count = 15310;
	#10 counter$count = 15311;
	#10 counter$count = 15312;
	#10 counter$count = 15313;
	#10 counter$count = 15314;
	#10 counter$count = 15315;
	#10 counter$count = 15316;
	#10 counter$count = 15317;
	#10 counter$count = 15318;
	#10 counter$count = 15319;
	#10 counter$count = 15320;
	#10 counter$count = 15321;
	#10 counter$count = 15322;
	#10 counter$count = 15323;
	#10 counter$count = 15324;
	#10 counter$count = 15325;
	#10 counter$count = 15326;
	#10 counter$count = 15327;
	#10 counter$count = 15328;
	#10 counter$count = 15329;
	#10 counter$count = 15330;
	#10 counter$count = 15331;
	#10 counter$count = 15332;
	#10 counter$count = 15333;
	#10 counter$count = 15334;
	#10 counter$count = 15335;
	#10 counter$count = 15336;
	#10 counter$count = 15337;
	#10 counter$count = 15338;
	#10 counter$count = 15339;
	#10 counter$count = 15340;
	#10 counter$count = 15341;
	#10 counter$count = 15342;
	#10 counter$count = 15343;
	#10 counter$count = 15344;
	#10 counter$count = 15345;
	#10 counter$count = 15346;
	#10 counter$count = 15347;
	#10 counter$count = 15348;
	#10 counter$count = 15349;
	#10 counter$count = 15350;
	#10 counter$count = 15351;
	#10 counter$count = 15352;
	#10 counter$count = 15353;
	#10 counter$count = 15354;
	#10 counter$count = 15355;
	#10 counter$count = 15356;
	#10 counter$count = 15357;
	#10 counter$count = 15358;
	#10 counter$count = 15359;
	#10 counter$count = 15360;
	#10 counter$count = 15361;
	#10 counter$count = 15362;
	#10 counter$count = 15363;
	#10 counter$count = 15364;
	#10 counter$count = 15365;
	#10 counter$count = 15366;
	#10 counter$count = 15367;
	#10 counter$count = 15368;
	#10 counter$count = 15369;
	#10 counter$count = 15370;
	#10 counter$count = 15371;
	#10 counter$count = 15372;
	#10 counter$count = 15373;
	#10 counter$count = 15374;
	#10 counter$count = 15375;
	#10 counter$count = 15376;
	#10 counter$count = 15377;
	#10 counter$count = 15378;
	#10 counter$count = 15379;
	#10 counter$count = 15380;
	#10 counter$count = 15381;
	#10 counter$count = 15382;
	#10 counter$count = 15383;
	#10 counter$count = 15384;
	#10 counter$count = 15385;
	#10 counter$count = 15386;
	#10 counter$count = 15387;
	#10 counter$count = 15388;
	#10 counter$count = 15389;
	#10 counter$count = 15390;
	#10 counter$count = 15391;
	#10 counter$count = 15392;
	#10 counter$count = 15393;
	#10 counter$count = 15394;
	#10 counter$count = 15395;
	#10 counter$count = 15396;
	#10 counter$count = 15397;
	#10 counter$count = 15398;
	#10 counter$count = 15399;
	#10 counter$count = 15400;
	#10 counter$count = 15401;
	#10 counter$count = 15402;
	#10 counter$count = 15403;
	#10 counter$count = 15404;
	#10 counter$count = 15405;
	#10 counter$count = 15406;
	#10 counter$count = 15407;
	#10 counter$count = 15408;
	#10 counter$count = 15409;
	#10 counter$count = 15410;
	#10 counter$count = 15411;
	#10 counter$count = 15412;
	#10 counter$count = 15413;
	#10 counter$count = 15414;
	#10 counter$count = 15415;
	#10 counter$count = 15416;
	#10 counter$count = 15417;
	#10 counter$count = 15418;
	#10 counter$count = 15419;
	#10 counter$count = 15420;
	#10 counter$count = 15421;
	#10 counter$count = 15422;
	#10 counter$count = 15423;
	#10 counter$count = 15424;
	#10 counter$count = 15425;
	#10 counter$count = 15426;
	#10 counter$count = 15427;
	#10 counter$count = 15428;
	#10 counter$count = 15429;
	#10 counter$count = 15430;
	#10 counter$count = 15431;
	#10 counter$count = 15432;
	#10 counter$count = 15433;
	#10 counter$count = 15434;
	#10 counter$count = 15435;
	#10 counter$count = 15436;
	#10 counter$count = 15437;
	#10 counter$count = 15438;
	#10 counter$count = 15439;
	#10 counter$count = 15440;
	#10 counter$count = 15441;
	#10 counter$count = 15442;
	#10 counter$count = 15443;
	#10 counter$count = 15444;
	#10 counter$count = 15445;
	#10 counter$count = 15446;
	#10 counter$count = 15447;
	#10 counter$count = 15448;
	#10 counter$count = 15449;
	#10 counter$count = 15450;
	#10 counter$count = 15451;
	#10 counter$count = 15452;
	#10 counter$count = 15453;
	#10 counter$count = 15454;
	#10 counter$count = 15455;
	#10 counter$count = 15456;
	#10 counter$count = 15457;
	#10 counter$count = 15458;
	#10 counter$count = 15459;
	#10 counter$count = 15460;
	#10 counter$count = 15461;
	#10 counter$count = 15462;
	#10 counter$count = 15463;
	#10 counter$count = 15464;
	#10 counter$count = 15465;
	#10 counter$count = 15466;
	#10 counter$count = 15467;
	#10 counter$count = 15468;
	#10 counter$count = 15469;
	#10 counter$count = 15470;
	#10 counter$count = 15471;
	#10 counter$count = 15472;
	#10 counter$count = 15473;
	#10 counter$count = 15474;
	#10 counter$count = 15475;
	#10 counter$count = 15476;
	#10 counter$count = 15477;
	#10 counter$count = 15478;
	#10 counter$count = 15479;
	#10 counter$count = 15480;
	#10 counter$count = 15481;
	#10 counter$count = 15482;
	#10 counter$count = 15483;
	#10 counter$count = 15484;
	#10 counter$count = 15485;
	#10 counter$count = 15486;
	#10 counter$count = 15487;
	#10 counter$count = 15488;
	#10 counter$count = 15489;
	#10 counter$count = 15490;
	#10 counter$count = 15491;
	#10 counter$count = 15492;
	#10 counter$count = 15493;
	#10 counter$count = 15494;
	#10 counter$count = 15495;
	#10 counter$count = 15496;
	#10 counter$count = 15497;
	#10 counter$count = 15498;
	#10 counter$count = 15499;
	#10 counter$count = 15500;
	#10 counter$count = 15501;
	#10 counter$count = 15502;
	#10 counter$count = 15503;
	#10 counter$count = 15504;
	#10 counter$count = 15505;
	#10 counter$count = 15506;
	#10 counter$count = 15507;
	#10 counter$count = 15508;
	#10 counter$count = 15509;
	#10 counter$count = 15510;
	#10 counter$count = 15511;
	#10 counter$count = 15512;
	#10 counter$count = 15513;
	#10 counter$count = 15514;
	#10 counter$count = 15515;
	#10 counter$count = 15516;
	#10 counter$count = 15517;
	#10 counter$count = 15518;
	#10 counter$count = 15519;
	#10 counter$count = 15520;
	#10 counter$count = 15521;
	#10 counter$count = 15522;
	#10 counter$count = 15523;
	#10 counter$count = 15524;
	#10 counter$count = 15525;
	#10 counter$count = 15526;
	#10 counter$count = 15527;
	#10 counter$count = 15528;
	#10 counter$count = 15529;
	#10 counter$count = 15530;
	#10 counter$count = 15531;
	#10 counter$count = 15532;
	#10 counter$count = 15533;
	#10 counter$count = 15534;
	#10 counter$count = 15535;
	#10 counter$count = 15536;
	#10 counter$count = 15537;
	#10 counter$count = 15538;
	#10 counter$count = 15539;
	#10 counter$count = 15540;
	#10 counter$count = 15541;
	#10 counter$count = 15542;
	#10 counter$count = 15543;
	#10 counter$count = 15544;
	#10 counter$count = 15545;
	#10 counter$count = 15546;
	#10 counter$count = 15547;
	#10 counter$count = 15548;
	#10 counter$count = 15549;
	#10 counter$count = 15550;
	#10 counter$count = 15551;
	#10 counter$count = 15552;
	#10 counter$count = 15553;
	#10 counter$count = 15554;
	#10 counter$count = 15555;
	#10 counter$count = 15556;
	#10 counter$count = 15557;
	#10 counter$count = 15558;
	#10 counter$count = 15559;
	#10 counter$count = 15560;
	#10 counter$count = 15561;
	#10 counter$count = 15562;
	#10 counter$count = 15563;
	#10 counter$count = 15564;
	#10 counter$count = 15565;
	#10 counter$count = 15566;
	#10 counter$count = 15567;
	#10 counter$count = 15568;
	#10 counter$count = 15569;
	#10 counter$count = 15570;
	#10 counter$count = 15571;
	#10 counter$count = 15572;
	#10 counter$count = 15573;
	#10 counter$count = 15574;
	#10 counter$count = 15575;
	#10 counter$count = 15576;
	#10 counter$count = 15577;
	#10 counter$count = 15578;
	#10 counter$count = 15579;
	#10 counter$count = 15580;
	#10 counter$count = 15581;
	#10 counter$count = 15582;
	#10 counter$count = 15583;
	#10 counter$count = 15584;
	#10 counter$count = 15585;
	#10 counter$count = 15586;
	#10 counter$count = 15587;
	#10 counter$count = 15588;
	#10 counter$count = 15589;
	#10 counter$count = 15590;
	#10 counter$count = 15591;
	#10 counter$count = 15592;
	#10 counter$count = 15593;
	#10 counter$count = 15594;
	#10 counter$count = 15595;
	#10 counter$count = 15596;
	#10 counter$count = 15597;
	#10 counter$count = 15598;
	#10 counter$count = 15599;
	#10 counter$count = 15600;
	#10 counter$count = 15601;
	#10 counter$count = 15602;
	#10 counter$count = 15603;
	#10 counter$count = 15604;
	#10 counter$count = 15605;
	#10 counter$count = 15606;
	#10 counter$count = 15607;
	#10 counter$count = 15608;
	#10 counter$count = 15609;
	#10 counter$count = 15610;
	#10 counter$count = 15611;
	#10 counter$count = 15612;
	#10 counter$count = 15613;
	#10 counter$count = 15614;
	#10 counter$count = 15615;
	#10 counter$count = 15616;
	#10 counter$count = 15617;
	#10 counter$count = 15618;
	#10 counter$count = 15619;
	#10 counter$count = 15620;
	#10 counter$count = 15621;
	#10 counter$count = 15622;
	#10 counter$count = 15623;
	#10 counter$count = 15624;
	#10 counter$count = 15625;
	#10 counter$count = 15626;
	#10 counter$count = 15627;
	#10 counter$count = 15628;
	#10 counter$count = 15629;
	#10 counter$count = 15630;
	#10 counter$count = 15631;
	#10 counter$count = 15632;
	#10 counter$count = 15633;
	#10 counter$count = 15634;
	#10 counter$count = 15635;
	#10 counter$count = 15636;
	#10 counter$count = 15637;
	#10 counter$count = 15638;
	#10 counter$count = 15639;
	#10 counter$count = 15640;
	#10 counter$count = 15641;
	#10 counter$count = 15642;
	#10 counter$count = 15643;
	#10 counter$count = 15644;
	#10 counter$count = 15645;
	#10 counter$count = 15646;
	#10 counter$count = 15647;
	#10 counter$count = 15648;
	#10 counter$count = 15649;
	#10 counter$count = 15650;
	#10 counter$count = 15651;
	#10 counter$count = 15652;
	#10 counter$count = 15653;
	#10 counter$count = 15654;
	#10 counter$count = 15655;
	#10 counter$count = 15656;
	#10 counter$count = 15657;
	#10 counter$count = 15658;
	#10 counter$count = 15659;
	#10 counter$count = 15660;
	#10 counter$count = 15661;
	#10 counter$count = 15662;
	#10 counter$count = 15663;
	#10 counter$count = 15664;
	#10 counter$count = 15665;
	#10 counter$count = 15666;
	#10 counter$count = 15667;
	#10 counter$count = 15668;
	#10 counter$count = 15669;
	#10 counter$count = 15670;
	#10 counter$count = 15671;
	#10 counter$count = 15672;
	#10 counter$count = 15673;
	#10 counter$count = 15674;
	#10 counter$count = 15675;
	#10 counter$count = 15676;
	#10 counter$count = 15677;
	#10 counter$count = 15678;
	#10 counter$count = 15679;
	#10 counter$count = 15680;
	#10 counter$count = 15681;
	#10 counter$count = 15682;
	#10 counter$count = 15683;
	#10 counter$count = 15684;
	#10 counter$count = 15685;
	#10 counter$count = 15686;
	#10 counter$count = 15687;
	#10 counter$count = 15688;
	#10 counter$count = 15689;
	#10 counter$count = 15690;
	#10 counter$count = 15691;
	#10 counter$count = 15692;
	#10 counter$count = 15693;
	#10 counter$count = 15694;
	#10 counter$count = 15695;
	#10 counter$count = 15696;
	#10 counter$count = 15697;
	#10 counter$count = 15698;
	#10 counter$count = 15699;
	#10 counter$count = 15700;
	#10 counter$count = 15701;
	#10 counter$count = 15702;
	#10 counter$count = 15703;
	#10 counter$count = 15704;
	#10 counter$count = 15705;
	#10 counter$count = 15706;
	#10 counter$count = 15707;
	#10 counter$count = 15708;
	#10 counter$count = 15709;
	#10 counter$count = 15710;
	#10 counter$count = 15711;
	#10 counter$count = 15712;
	#10 counter$count = 15713;
	#10 counter$count = 15714;
	#10 counter$count = 15715;
	#10 counter$count = 15716;
	#10 counter$count = 15717;
	#10 counter$count = 15718;
	#10 counter$count = 15719;
	#10 counter$count = 15720;
	#10 counter$count = 15721;
	#10 counter$count = 15722;
	#10 counter$count = 15723;
	#10 counter$count = 15724;
	#10 counter$count = 15725;
	#10 counter$count = 15726;
	#10 counter$count = 15727;
	#10 counter$count = 15728;
	#10 counter$count = 15729;
	#10 counter$count = 15730;
	#10 counter$count = 15731;
	#10 counter$count = 15732;
	#10 counter$count = 15733;
	#10 counter$count = 15734;
	#10 counter$count = 15735;
	#10 counter$count = 15736;
	#10 counter$count = 15737;
	#10 counter$count = 15738;
	#10 counter$count = 15739;
	#10 counter$count = 15740;
	#10 counter$count = 15741;
	#10 counter$count = 15742;
	#10 counter$count = 15743;
	#10 counter$count = 15744;
	#10 counter$count = 15745;
	#10 counter$count = 15746;
	#10 counter$count = 15747;
	#10 counter$count = 15748;
	#10 counter$count = 15749;
	#10 counter$count = 15750;
	#10 counter$count = 15751;
	#10 counter$count = 15752;
	#10 counter$count = 15753;
	#10 counter$count = 15754;
	#10 counter$count = 15755;
	#10 counter$count = 15756;
	#10 counter$count = 15757;
	#10 counter$count = 15758;
	#10 counter$count = 15759;
	#10 counter$count = 15760;
	#10 counter$count = 15761;
	#10 counter$count = 15762;
	#10 counter$count = 15763;
	#10 counter$count = 15764;
	#10 counter$count = 15765;
	#10 counter$count = 15766;
	#10 counter$count = 15767;
	#10 counter$count = 15768;
	#10 counter$count = 15769;
	#10 counter$count = 15770;
	#10 counter$count = 15771;
	#10 counter$count = 15772;
	#10 counter$count = 15773;
	#10 counter$count = 15774;
	#10 counter$count = 15775;
	#10 counter$count = 15776;
	#10 counter$count = 15777;
	#10 counter$count = 15778;
	#10 counter$count = 15779;
	#10 counter$count = 15780;
	#10 counter$count = 15781;
	#10 counter$count = 15782;
	#10 counter$count = 15783;
	#10 counter$count = 15784;
	#10 counter$count = 15785;
	#10 counter$count = 15786;
	#10 counter$count = 15787;
	#10 counter$count = 15788;
	#10 counter$count = 15789;
	#10 counter$count = 15790;
	#10 counter$count = 15791;
	#10 counter$count = 15792;
	#10 counter$count = 15793;
	#10 counter$count = 15794;
	#10 counter$count = 15795;
	#10 counter$count = 15796;
	#10 counter$count = 15797;
	#10 counter$count = 15798;
	#10 counter$count = 15799;
	#10 counter$count = 15800;
	#10 counter$count = 15801;
	#10 counter$count = 15802;
	#10 counter$count = 15803;
	#10 counter$count = 15804;
	#10 counter$count = 15805;
	#10 counter$count = 15806;
	#10 counter$count = 15807;
	#10 counter$count = 15808;
	#10 counter$count = 15809;
	#10 counter$count = 15810;
	#10 counter$count = 15811;
	#10 counter$count = 15812;
	#10 counter$count = 15813;
	#10 counter$count = 15814;
	#10 counter$count = 15815;
	#10 counter$count = 15816;
	#10 counter$count = 15817;
	#10 counter$count = 15818;
	#10 counter$count = 15819;
	#10 counter$count = 15820;
	#10 counter$count = 15821;
	#10 counter$count = 15822;
	#10 counter$count = 15823;
	#10 counter$count = 15824;
	#10 counter$count = 15825;
	#10 counter$count = 15826;
	#10 counter$count = 15827;
	#10 counter$count = 15828;
	#10 counter$count = 15829;
	#10 counter$count = 15830;
	#10 counter$count = 15831;
	#10 counter$count = 15832;
	#10 counter$count = 15833;
	#10 counter$count = 15834;
	#10 counter$count = 15835;
	#10 counter$count = 15836;
	#10 counter$count = 15837;
	#10 counter$count = 15838;
	#10 counter$count = 15839;
	#10 counter$count = 15840;
	#10 counter$count = 15841;
	#10 counter$count = 15842;
	#10 counter$count = 15843;
	#10 counter$count = 15844;
	#10 counter$count = 15845;
	#10 counter$count = 15846;
	#10 counter$count = 15847;
	#10 counter$count = 15848;
	#10 counter$count = 15849;
	#10 counter$count = 15850;
	#10 counter$count = 15851;
	#10 counter$count = 15852;
	#10 counter$count = 15853;
	#10 counter$count = 15854;
	#10 counter$count = 15855;
	#10 counter$count = 15856;
	#10 counter$count = 15857;
	#10 counter$count = 15858;
	#10 counter$count = 15859;
	#10 counter$count = 15860;
	#10 counter$count = 15861;
	#10 counter$count = 15862;
	#10 counter$count = 15863;
	#10 counter$count = 15864;
	#10 counter$count = 15865;
	#10 counter$count = 15866;
	#10 counter$count = 15867;
	#10 counter$count = 15868;
	#10 counter$count = 15869;
	#10 counter$count = 15870;
	#10 counter$count = 15871;
	#10 counter$count = 15872;
	#10 counter$count = 15873;
	#10 counter$count = 15874;
	#10 counter$count = 15875;
	#10 counter$count = 15876;
	#10 counter$count = 15877;
	#10 counter$count = 15878;
	#10 counter$count = 15879;
	#10 counter$count = 15880;
	#10 counter$count = 15881;
	#10 counter$count = 15882;
	#10 counter$count = 15883;
	#10 counter$count = 15884;
	#10 counter$count = 15885;
	#10 counter$count = 15886;
	#10 counter$count = 15887;
	#10 counter$count = 15888;
	#10 counter$count = 15889;
	#10 counter$count = 15890;
	#10 counter$count = 15891;
	#10 counter$count = 15892;
	#10 counter$count = 15893;
	#10 counter$count = 15894;
	#10 counter$count = 15895;
	#10 counter$count = 15896;
	#10 counter$count = 15897;
	#10 counter$count = 15898;
	#10 counter$count = 15899;
	#10 counter$count = 15900;
	#10 counter$count = 15901;
	#10 counter$count = 15902;
	#10 counter$count = 15903;
	#10 counter$count = 15904;
	#10 counter$count = 15905;
	#10 counter$count = 15906;
	#10 counter$count = 15907;
	#10 counter$count = 15908;
	#10 counter$count = 15909;
	#10 counter$count = 15910;
	#10 counter$count = 15911;
	#10 counter$count = 15912;
	#10 counter$count = 15913;
	#10 counter$count = 15914;
	#10 counter$count = 15915;
	#10 counter$count = 15916;
	#10 counter$count = 15917;
	#10 counter$count = 15918;
	#10 counter$count = 15919;
	#10 counter$count = 15920;
	#10 counter$count = 15921;
	#10 counter$count = 15922;
	#10 counter$count = 15923;
	#10 counter$count = 15924;
	#10 counter$count = 15925;
	#10 counter$count = 15926;
	#10 counter$count = 15927;
	#10 counter$count = 15928;
	#10 counter$count = 15929;
	#10 counter$count = 15930;
	#10 counter$count = 15931;
	#10 counter$count = 15932;
	#10 counter$count = 15933;
	#10 counter$count = 15934;
	#10 counter$count = 15935;
	#10 counter$count = 15936;
	#10 counter$count = 15937;
	#10 counter$count = 15938;
	#10 counter$count = 15939;
	#10 counter$count = 15940;
	#10 counter$count = 15941;
	#10 counter$count = 15942;
	#10 counter$count = 15943;
	#10 counter$count = 15944;
	#10 counter$count = 15945;
	#10 counter$count = 15946;
	#10 counter$count = 15947;
	#10 counter$count = 15948;
	#10 counter$count = 15949;
	#10 counter$count = 15950;
	#10 counter$count = 15951;
	#10 counter$count = 15952;
	#10 counter$count = 15953;
	#10 counter$count = 15954;
	#10 counter$count = 15955;
	#10 counter$count = 15956;
	#10 counter$count = 15957;
	#10 counter$count = 15958;
	#10 counter$count = 15959;
	#10 counter$count = 15960;
	#10 counter$count = 15961;
	#10 counter$count = 15962;
	#10 counter$count = 15963;
	#10 counter$count = 15964;
	#10 counter$count = 15965;
	#10 counter$count = 15966;
	#10 counter$count = 15967;
	#10 counter$count = 15968;
	#10 counter$count = 15969;
	#10 counter$count = 15970;
	#10 counter$count = 15971;
	#10 counter$count = 15972;
	#10 counter$count = 15973;
	#10 counter$count = 15974;
	#10 counter$count = 15975;
	#10 counter$count = 15976;
	#10 counter$count = 15977;
	#10 counter$count = 15978;
	#10 counter$count = 15979;
	#10 counter$count = 15980;
	#10 counter$count = 15981;
	#10 counter$count = 15982;
	#10 counter$count = 15983;
	#10 counter$count = 15984;
	#10 counter$count = 15985;
	#10 counter$count = 15986;
	#10 counter$count = 15987;
	#10 counter$count = 15988;
	#10 counter$count = 15989;
	#10 counter$count = 15990;
	#10 counter$count = 15991;
	#10 counter$count = 15992;
	#10 counter$count = 15993;
	#10 counter$count = 15994;
	#10 counter$count = 15995;
	#10 counter$count = 15996;
	#10 counter$count = 15997;
	#10 counter$count = 15998;
	#10 counter$count = 15999;
	#10 counter$count = 16000;
	#10 counter$count = 16001;
	#10 counter$count = 16002;
	#10 counter$count = 16003;
	#10 counter$count = 16004;
	#10 counter$count = 16005;
	#10 counter$count = 16006;
	#10 counter$count = 16007;
	#10 counter$count = 16008;
	#10 counter$count = 16009;
	#10 counter$count = 16010;
	#10 counter$count = 16011;
	#10 counter$count = 16012;
	#10 counter$count = 16013;
	#10 counter$count = 16014;
	#10 counter$count = 16015;
	#10 counter$count = 16016;
	#10 counter$count = 16017;
	#10 counter$count = 16018;
	#10 counter$count = 16019;
	#10 counter$count = 16020;
	#10 counter$count = 16021;
	#10 counter$count = 16022;
	#10 counter$count = 16023;
	#10 counter$count = 16024;
	#10 counter$count = 16025;
	#10 counter$count = 16026;
	#10 counter$count = 16027;
	#10 counter$count = 16028;
	#10 counter$count = 16029;
	#10 counter$count = 16030;
	#10 counter$count = 16031;
	#10 counter$count = 16032;
	#10 counter$count = 16033;
	#10 counter$count = 16034;
	#10 counter$count = 16035;
	#10 counter$count = 16036;
	#10 counter$count = 16037;
	#10 counter$count = 16038;
	#10 counter$count = 16039;
	#10 counter$count = 16040;
	#10 counter$count = 16041;
	#10 counter$count = 16042;
	#10 counter$count = 16043;
	#10 counter$count = 16044;
	#10 counter$count = 16045;
	#10 counter$count = 16046;
	#10 counter$count = 16047;
	#10 counter$count = 16048;
	#10 counter$count = 16049;
	#10 counter$count = 16050;
	#10 counter$count = 16051;
	#10 counter$count = 16052;
	#10 counter$count = 16053;
	#10 counter$count = 16054;
	#10 counter$count = 16055;
	#10 counter$count = 16056;
	#10 counter$count = 16057;
	#10 counter$count = 16058;
	#10 counter$count = 16059;
	#10 counter$count = 16060;
	#10 counter$count = 16061;
	#10 counter$count = 16062;
	#10 counter$count = 16063;
	#10 counter$count = 16064;
	#10 counter$count = 16065;
	#10 counter$count = 16066;
	#10 counter$count = 16067;
	#10 counter$count = 16068;
	#10 counter$count = 16069;
	#10 counter$count = 16070;
	#10 counter$count = 16071;
	#10 counter$count = 16072;
	#10 counter$count = 16073;
	#10 counter$count = 16074;
	#10 counter$count = 16075;
	#10 counter$count = 16076;
	#10 counter$count = 16077;
	#10 counter$count = 16078;
	#10 counter$count = 16079;
	#10 counter$count = 16080;
	#10 counter$count = 16081;
	#10 counter$count = 16082;
	#10 counter$count = 16083;
	#10 counter$count = 16084;
	#10 counter$count = 16085;
	#10 counter$count = 16086;
	#10 counter$count = 16087;
	#10 counter$count = 16088;
	#10 counter$count = 16089;
	#10 counter$count = 16090;
	#10 counter$count = 16091;
	#10 counter$count = 16092;
	#10 counter$count = 16093;
	#10 counter$count = 16094;
	#10 counter$count = 16095;
	#10 counter$count = 16096;
	#10 counter$count = 16097;
	#10 counter$count = 16098;
	#10 counter$count = 16099;
	#10 counter$count = 16100;
	#10 counter$count = 16101;
	#10 counter$count = 16102;
	#10 counter$count = 16103;
	#10 counter$count = 16104;
	#10 counter$count = 16105;
	#10 counter$count = 16106;
	#10 counter$count = 16107;
	#10 counter$count = 16108;
	#10 counter$count = 16109;
	#10 counter$count = 16110;
	#10 counter$count = 16111;
	#10 counter$count = 16112;
	#10 counter$count = 16113;
	#10 counter$count = 16114;
	#10 counter$count = 16115;
	#10 counter$count = 16116;
	#10 counter$count = 16117;
	#10 counter$count = 16118;
	#10 counter$count = 16119;
	#10 counter$count = 16120;
	#10 counter$count = 16121;
	#10 counter$count = 16122;
	#10 counter$count = 16123;
	#10 counter$count = 16124;
	#10 counter$count = 16125;
	#10 counter$count = 16126;
	#10 counter$count = 16127;
	#10 counter$count = 16128;
	#10 counter$count = 16129;
	#10 counter$count = 16130;
	#10 counter$count = 16131;
	#10 counter$count = 16132;
	#10 counter$count = 16133;
	#10 counter$count = 16134;
	#10 counter$count = 16135;
	#10 counter$count = 16136;
	#10 counter$count = 16137;
	#10 counter$count = 16138;
	#10 counter$count = 16139;
	#10 counter$count = 16140;
	#10 counter$count = 16141;
	#10 counter$count = 16142;
	#10 counter$count = 16143;
	#10 counter$count = 16144;
	#10 counter$count = 16145;
	#10 counter$count = 16146;
	#10 counter$count = 16147;
	#10 counter$count = 16148;
	#10 counter$count = 16149;
	#10 counter$count = 16150;
	#10 counter$count = 16151;
	#10 counter$count = 16152;
	#10 counter$count = 16153;
	#10 counter$count = 16154;
	#10 counter$count = 16155;
	#10 counter$count = 16156;
	#10 counter$count = 16157;
	#10 counter$count = 16158;
	#10 counter$count = 16159;
	#10 counter$count = 16160;
	#10 counter$count = 16161;
	#10 counter$count = 16162;
	#10 counter$count = 16163;
	#10 counter$count = 16164;
	#10 counter$count = 16165;
	#10 counter$count = 16166;
	#10 counter$count = 16167;
	#10 counter$count = 16168;
	#10 counter$count = 16169;
	#10 counter$count = 16170;
	#10 counter$count = 16171;
	#10 counter$count = 16172;
	#10 counter$count = 16173;
	#10 counter$count = 16174;
	#10 counter$count = 16175;
	#10 counter$count = 16176;
	#10 counter$count = 16177;
	#10 counter$count = 16178;
	#10 counter$count = 16179;
	#10 counter$count = 16180;
	#10 counter$count = 16181;
	#10 counter$count = 16182;
	#10 counter$count = 16183;
	#10 counter$count = 16184;
	#10 counter$count = 16185;
	#10 counter$count = 16186;
	#10 counter$count = 16187;
	#10 counter$count = 16188;
	#10 counter$count = 16189;
	#10 counter$count = 16190;
	#10 counter$count = 16191;
	#10 counter$count = 16192;
	#10 counter$count = 16193;
	#10 counter$count = 16194;
	#10 counter$count = 16195;
	#10 counter$count = 16196;
	#10 counter$count = 16197;
	#10 counter$count = 16198;
	#10 counter$count = 16199;
	#10 counter$count = 16200;
	#10 counter$count = 16201;
	#10 counter$count = 16202;
	#10 counter$count = 16203;
	#10 counter$count = 16204;
	#10 counter$count = 16205;
	#10 counter$count = 16206;
	#10 counter$count = 16207;
	#10 counter$count = 16208;
	#10 counter$count = 16209;
	#10 counter$count = 16210;
	#10 counter$count = 16211;
	#10 counter$count = 16212;
	#10 counter$count = 16213;
	#10 counter$count = 16214;
	#10 counter$count = 16215;
	#10 counter$count = 16216;
	#10 counter$count = 16217;
	#10 counter$count = 16218;
	#10 counter$count = 16219;
	#10 counter$count = 16220;
	#10 counter$count = 16221;
	#10 counter$count = 16222;
	#10 counter$count = 16223;
	#10 counter$count = 16224;
	#10 counter$count = 16225;
	#10 counter$count = 16226;
	#10 counter$count = 16227;
	#10 counter$count = 16228;
	#10 counter$count = 16229;
	#10 counter$count = 16230;
	#10 counter$count = 16231;
	#10 counter$count = 16232;
	#10 counter$count = 16233;
	#10 counter$count = 16234;
	#10 counter$count = 16235;
	#10 counter$count = 16236;
	#10 counter$count = 16237;
	#10 counter$count = 16238;
	#10 counter$count = 16239;
	#10 counter$count = 16240;
	#10 counter$count = 16241;
	#10 counter$count = 16242;
	#10 counter$count = 16243;
	#10 counter$count = 16244;
	#10 counter$count = 16245;
	#10 counter$count = 16246;
	#10 counter$count = 16247;
	#10 counter$count = 16248;
	#10 counter$count = 16249;
	#10 counter$count = 16250;
	#10 counter$count = 16251;
	#10 counter$count = 16252;
	#10 counter$count = 16253;
	#10 counter$count = 16254;
	#10 counter$count = 16255;
	#10 counter$count = 16256;
	#10 counter$count = 16257;
	#10 counter$count = 16258;
	#10 counter$count = 16259;
	#10 counter$count = 16260;
	#10 counter$count = 16261;
	#10 counter$count = 16262;
	#10 counter$count = 16263;
	#10 counter$count = 16264;
	#10 counter$count = 16265;
	#10 counter$count = 16266;
	#10 counter$count = 16267;
	#10 counter$count = 16268;
	#10 counter$count = 16269;
	#10 counter$count = 16270;
	#10 counter$count = 16271;
	#10 counter$count = 16272;
	#10 counter$count = 16273;
	#10 counter$count = 16274;
	#10 counter$count = 16275;
	#10 counter$count = 16276;
	#10 counter$count = 16277;
	#10 counter$count = 16278;
	#10 counter$count = 16279;
	#10 counter$count = 16280;
	#10 counter$count = 16281;
	#10 counter$count = 16282;
	#10 counter$count = 16283;
	#10 counter$count = 16284;
	#10 counter$count = 16285;
	#10 counter$count = 16286;
	#10 counter$count = 16287;
	#10 counter$count = 16288;
	#10 counter$count = 16289;
	#10 counter$count = 16290;
	#10 counter$count = 16291;
	#10 counter$count = 16292;
	#10 counter$count = 16293;
	#10 counter$count = 16294;
	#10 counter$count = 16295;
	#10 counter$count = 16296;
	#10 counter$count = 16297;
	#10 counter$count = 16298;
	#10 counter$count = 16299;
	#10 counter$count = 16300;
	#10 counter$count = 16301;
	#10 counter$count = 16302;
	#10 counter$count = 16303;
	#10 counter$count = 16304;
	#10 counter$count = 16305;
	#10 counter$count = 16306;
	#10 counter$count = 16307;
	#10 counter$count = 16308;
	#10 counter$count = 16309;
	#10 counter$count = 16310;
	#10 counter$count = 16311;
	#10 counter$count = 16312;
	#10 counter$count = 16313;
	#10 counter$count = 16314;
	#10 counter$count = 16315;
	#10 counter$count = 16316;
	#10 counter$count = 16317;
	#10 counter$count = 16318;
	#10 counter$count = 16319;
	#10 counter$count = 16320;
	#10 counter$count = 16321;
	#10 counter$count = 16322;
	#10 counter$count = 16323;
	#10 counter$count = 16324;
	#10 counter$count = 16325;
	#10 counter$count = 16326;
	#10 counter$count = 16327;
	#10 counter$count = 16328;
	#10 counter$count = 16329;
	#10 counter$count = 16330;
	#10 counter$count = 16331;
	#10 counter$count = 16332;
	#10 counter$count = 16333;
	#10 counter$count = 16334;
	#10 counter$count = 16335;
	#10 counter$count = 16336;
	#10 counter$count = 16337;
	#10 counter$count = 16338;
	#10 counter$count = 16339;
	#10 counter$count = 16340;
	#10 counter$count = 16341;
	#10 counter$count = 16342;
	#10 counter$count = 16343;
	#10 counter$count = 16344;
	#10 counter$count = 16345;
	#10 counter$count = 16346;
	#10 counter$count = 16347;
	#10 counter$count = 16348;
	#10 counter$count = 16349;
	#10 counter$count = 16350;
	#10 counter$count = 16351;
	#10 counter$count = 16352;
	#10 counter$count = 16353;
	#10 counter$count = 16354;
	#10 counter$count = 16355;
	#10 counter$count = 16356;
	#10 counter$count = 16357;
	#10 counter$count = 16358;
	#10 counter$count = 16359;
	#10 counter$count = 16360;
	#10 counter$count = 16361;
	#10 counter$count = 16362;
	#10 counter$count = 16363;
	#10 counter$count = 16364;
	#10 counter$count = 16365;
	#10 counter$count = 16366;
	#10 counter$count = 16367;
	#10 counter$count = 16368;
	#10 counter$count = 16369;
	#10 counter$count = 16370;
	#10 counter$count = 16371;
	#10 counter$count = 16372;
	#10 counter$count = 16373;
	#10 counter$count = 16374;
	#10 counter$count = 16375;
	#10 counter$count = 16376;
	#10 counter$count = 16377;
	#10 counter$count = 16378;
	#10 counter$count = 16379;
	#10 counter$count = 16380;
	#10 counter$count = 16381;
	#10 counter$count = 16382;
	#10 counter$count = 16383;
	#10 counter$count = 16384;
	#10 counter$count = 16385;
	#10 counter$count = 16386;
	#10 counter$count = 16387;
	#10 counter$count = 16388;
	#10 counter$count = 16389;
	#10 counter$count = 16390;
	#10 counter$count = 16391;
	#10 counter$count = 16392;
	#10 counter$count = 16393;
	#10 counter$count = 16394;
	#10 counter$count = 16395;
	#10 counter$count = 16396;
	#10 counter$count = 16397;
	#10 counter$count = 16398;
	#10 counter$count = 16399;
	#10 counter$count = 16400;
	#10 counter$count = 16401;
	#10 counter$count = 16402;
	#10 counter$count = 16403;
	#10 counter$count = 16404;
	#10 counter$count = 16405;
	#10 counter$count = 16406;
	#10 counter$count = 16407;
	#10 counter$count = 16408;
	#10 counter$count = 16409;
	#10 counter$count = 16410;
	#10 counter$count = 16411;
	#10 counter$count = 16412;
	#10 counter$count = 16413;
	#10 counter$count = 16414;
	#10 counter$count = 16415;
	#10 counter$count = 16416;
	#10 counter$count = 16417;
	#10 counter$count = 16418;
	#10 counter$count = 16419;
	#10 counter$count = 16420;
	#10 counter$count = 16421;
	#10 counter$count = 16422;
	#10 counter$count = 16423;
	#10 counter$count = 16424;
	#10 counter$count = 16425;
	#10 counter$count = 16426;
	#10 counter$count = 16427;
	#10 counter$count = 16428;
	#10 counter$count = 16429;
	#10 counter$count = 16430;
	#10 counter$count = 16431;
	#10 counter$count = 16432;
	#10 counter$count = 16433;
	#10 counter$count = 16434;
	#10 counter$count = 16435;
	#10 counter$count = 16436;
	#10 counter$count = 16437;
	#10 counter$count = 16438;
	#10 counter$count = 16439;
	#10 counter$count = 16440;
	#10 counter$count = 16441;
	#10 counter$count = 16442;
	#10 counter$count = 16443;
	#10 counter$count = 16444;
	#10 counter$count = 16445;
	#10 counter$count = 16446;
	#10 counter$count = 16447;
	#10 counter$count = 16448;
	#10 counter$count = 16449;
	#10 counter$count = 16450;
	#10 counter$count = 16451;
	#10 counter$count = 16452;
	#10 counter$count = 16453;
	#10 counter$count = 16454;
	#10 counter$count = 16455;
	#10 counter$count = 16456;
	#10 counter$count = 16457;
	#10 counter$count = 16458;
	#10 counter$count = 16459;
	#10 counter$count = 16460;
	#10 counter$count = 16461;
	#10 counter$count = 16462;
	#10 counter$count = 16463;
	#10 counter$count = 16464;
	#10 counter$count = 16465;
	#10 counter$count = 16466;
	#10 counter$count = 16467;
	#10 counter$count = 16468;
	#10 counter$count = 16469;
	#10 counter$count = 16470;
	#10 counter$count = 16471;
	#10 counter$count = 16472;
	#10 counter$count = 16473;
	#10 counter$count = 16474;
	#10 counter$count = 16475;
	#10 counter$count = 16476;
	#10 counter$count = 16477;
	#10 counter$count = 16478;
	#10 counter$count = 16479;
	#10 counter$count = 16480;
	#10 counter$count = 16481;
	#10 counter$count = 16482;
	#10 counter$count = 16483;
	#10 counter$count = 16484;
	#10 counter$count = 16485;
	#10 counter$count = 16486;
	#10 counter$count = 16487;
	#10 counter$count = 16488;
	#10 counter$count = 16489;
	#10 counter$count = 16490;
	#10 counter$count = 16491;
	#10 counter$count = 16492;
	#10 counter$count = 16493;
	#10 counter$count = 16494;
	#10 counter$count = 16495;
	#10 counter$count = 16496;
	#10 counter$count = 16497;
	#10 counter$count = 16498;
	#10 counter$count = 16499;
	#10 counter$count = 16500;
	#10 counter$count = 16501;
	#10 counter$count = 16502;
	#10 counter$count = 16503;
	#10 counter$count = 16504;
	#10 counter$count = 16505;
	#10 counter$count = 16506;
	#10 counter$count = 16507;
	#10 counter$count = 16508;
	#10 counter$count = 16509;
	#10 counter$count = 16510;
	#10 counter$count = 16511;
	#10 counter$count = 16512;
	#10 counter$count = 16513;
	#10 counter$count = 16514;
	#10 counter$count = 16515;
	#10 counter$count = 16516;
	#10 counter$count = 16517;
	#10 counter$count = 16518;
	#10 counter$count = 16519;
	#10 counter$count = 16520;
	#10 counter$count = 16521;
	#10 counter$count = 16522;
	#10 counter$count = 16523;
	#10 counter$count = 16524;
	#10 counter$count = 16525;
	#10 counter$count = 16526;
	#10 counter$count = 16527;
	#10 counter$count = 16528;
	#10 counter$count = 16529;
	#10 counter$count = 16530;
	#10 counter$count = 16531;
	#10 counter$count = 16532;
	#10 counter$count = 16533;
	#10 counter$count = 16534;
	#10 counter$count = 16535;
	#10 counter$count = 16536;
	#10 counter$count = 16537;
	#10 counter$count = 16538;
	#10 counter$count = 16539;
	#10 counter$count = 16540;
	#10 counter$count = 16541;
	#10 counter$count = 16542;
	#10 counter$count = 16543;
	#10 counter$count = 16544;
	#10 counter$count = 16545;
	#10 counter$count = 16546;
	#10 counter$count = 16547;
	#10 counter$count = 16548;
	#10 counter$count = 16549;
	#10 counter$count = 16550;
	#10 counter$count = 16551;
	#10 counter$count = 16552;
	#10 counter$count = 16553;
	#10 counter$count = 16554;
	#10 counter$count = 16555;
	#10 counter$count = 16556;
	#10 counter$count = 16557;
	#10 counter$count = 16558;
	#10 counter$count = 16559;
	#10 counter$count = 16560;
	#10 counter$count = 16561;
	#10 counter$count = 16562;
	#10 counter$count = 16563;
	#10 counter$count = 16564;
	#10 counter$count = 16565;
	#10 counter$count = 16566;
	#10 counter$count = 16567;
	#10 counter$count = 16568;
	#10 counter$count = 16569;
	#10 counter$count = 16570;
	#10 counter$count = 16571;
	#10 counter$count = 16572;
	#10 counter$count = 16573;
	#10 counter$count = 16574;
	#10 counter$count = 16575;
	#10 counter$count = 16576;
	#10 counter$count = 16577;
	#10 counter$count = 16578;
	#10 counter$count = 16579;
	#10 counter$count = 16580;
	#10 counter$count = 16581;
	#10 counter$count = 16582;
	#10 counter$count = 16583;
	#10 counter$count = 16584;
	#10 counter$count = 16585;
	#10 counter$count = 16586;
	#10 counter$count = 16587;
	#10 counter$count = 16588;
	#10 counter$count = 16589;
	#10 counter$count = 16590;
	#10 counter$count = 16591;
	#10 counter$count = 16592;
	#10 counter$count = 16593;
	#10 counter$count = 16594;
	#10 counter$count = 16595;
	#10 counter$count = 16596;
	#10 counter$count = 16597;
	#10 counter$count = 16598;
	#10 counter$count = 16599;
	#10 counter$count = 16600;
	#10 counter$count = 16601;
	#10 counter$count = 16602;
	#10 counter$count = 16603;
	#10 counter$count = 16604;
	#10 counter$count = 16605;
	#10 counter$count = 16606;
	#10 counter$count = 16607;
	#10 counter$count = 16608;
	#10 counter$count = 16609;
	#10 counter$count = 16610;
	#10 counter$count = 16611;
	#10 counter$count = 16612;
	#10 counter$count = 16613;
	#10 counter$count = 16614;
	#10 counter$count = 16615;
	#10 counter$count = 16616;
	#10 counter$count = 16617;
	#10 counter$count = 16618;
	#10 counter$count = 16619;
	#10 counter$count = 16620;
	#10 counter$count = 16621;
	#10 counter$count = 16622;
	#10 counter$count = 16623;
	#10 counter$count = 16624;
	#10 counter$count = 16625;
	#10 counter$count = 16626;
	#10 counter$count = 16627;
	#10 counter$count = 16628;
	#10 counter$count = 16629;
	#10 counter$count = 16630;
	#10 counter$count = 16631;
	#10 counter$count = 16632;
	#10 counter$count = 16633;
	#10 counter$count = 16634;
	#10 counter$count = 16635;
	#10 counter$count = 16636;
	#10 counter$count = 16637;
	#10 counter$count = 16638;
	#10 counter$count = 16639;
	#10 counter$count = 16640;
	#10 counter$count = 16641;
	#10 counter$count = 16642;
	#10 counter$count = 16643;
	#10 counter$count = 16644;
	#10 counter$count = 16645;
	#10 counter$count = 16646;
	#10 counter$count = 16647;
	#10 counter$count = 16648;
	#10 counter$count = 16649;
	#10 counter$count = 16650;
	#10 counter$count = 16651;
	#10 counter$count = 16652;
	#10 counter$count = 16653;
	#10 counter$count = 16654;
	#10 counter$count = 16655;
	#10 counter$count = 16656;
	#10 counter$count = 16657;
	#10 counter$count = 16658;
	#10 counter$count = 16659;
	#10 counter$count = 16660;
	#10 counter$count = 16661;
	#10 counter$count = 16662;
	#10 counter$count = 16663;
	#10 counter$count = 16664;
	#10 counter$count = 16665;
	#10 counter$count = 16666;
	#10 counter$count = 16667;
	#10 counter$count = 16668;
	#10 counter$count = 16669;
	#10 counter$count = 16670;
	#10 counter$count = 16671;
	#10 counter$count = 16672;
	#10 counter$count = 16673;
	#10 counter$count = 16674;
	#10 counter$count = 16675;
	#10 counter$count = 16676;
	#10 counter$count = 16677;
	#10 counter$count = 16678;
	#10 counter$count = 16679;
	#10 counter$count = 16680;
	#10 counter$count = 16681;
	#10 counter$count = 16682;
	#10 counter$count = 16683;
	#10 counter$count = 16684;
	#10 counter$count = 16685;
	#10 counter$count = 16686;
	#10 counter$count = 16687;
	#10 counter$count = 16688;
	#10 counter$count = 16689;
	#10 counter$count = 16690;
	#10 counter$count = 16691;
	#10 counter$count = 16692;
	#10 counter$count = 16693;
	#10 counter$count = 16694;
	#10 counter$count = 16695;
	#10 counter$count = 16696;
	#10 counter$count = 16697;
	#10 counter$count = 16698;
	#10 counter$count = 16699;
	#10 counter$count = 16700;
	#10 counter$count = 16701;
	#10 counter$count = 16702;
	#10 counter$count = 16703;
	#10 counter$count = 16704;
	#10 counter$count = 16705;
	#10 counter$count = 16706;
	#10 counter$count = 16707;
	#10 counter$count = 16708;
	#10 counter$count = 16709;
	#10 counter$count = 16710;
	#10 counter$count = 16711;
	#10 counter$count = 16712;
	#10 counter$count = 16713;
	#10 counter$count = 16714;
	#10 counter$count = 16715;
	#10 counter$count = 16716;
	#10 counter$count = 16717;
	#10 counter$count = 16718;
	#10 counter$count = 16719;
	#10 counter$count = 16720;
	#10 counter$count = 16721;
	#10 counter$count = 16722;
	#10 counter$count = 16723;
	#10 counter$count = 16724;
	#10 counter$count = 16725;
	#10 counter$count = 16726;
	#10 counter$count = 16727;
	#10 counter$count = 16728;
	#10 counter$count = 16729;
	#10 counter$count = 16730;
	#10 counter$count = 16731;
	#10 counter$count = 16732;
	#10 counter$count = 16733;
	#10 counter$count = 16734;
	#10 counter$count = 16735;
	#10 counter$count = 16736;
	#10 counter$count = 16737;
	#10 counter$count = 16738;
	#10 counter$count = 16739;
	#10 counter$count = 16740;
	#10 counter$count = 16741;
	#10 counter$count = 16742;
	#10 counter$count = 16743;
	#10 counter$count = 16744;
	#10 counter$count = 16745;
	#10 counter$count = 16746;
	#10 counter$count = 16747;
	#10 counter$count = 16748;
	#10 counter$count = 16749;
	#10 counter$count = 16750;
	#10 counter$count = 16751;
	#10 counter$count = 16752;
	#10 counter$count = 16753;
	#10 counter$count = 16754;
	#10 counter$count = 16755;
	#10 counter$count = 16756;
	#10 counter$count = 16757;
	#10 counter$count = 16758;
	#10 counter$count = 16759;
	#10 counter$count = 16760;
	#10 counter$count = 16761;
	#10 counter$count = 16762;
	#10 counter$count = 16763;
	#10 counter$count = 16764;
	#10 counter$count = 16765;
	#10 counter$count = 16766;
	#10 counter$count = 16767;
	#10 counter$count = 16768;
	#10 counter$count = 16769;
	#10 counter$count = 16770;
	#10 counter$count = 16771;
	#10 counter$count = 16772;
	#10 counter$count = 16773;
	#10 counter$count = 16774;
	#10 counter$count = 16775;
	#10 counter$count = 16776;
	#10 counter$count = 16777;
	#10 counter$count = 16778;
	#10 counter$count = 16779;
	#10 counter$count = 16780;
	#10 counter$count = 16781;
	#10 counter$count = 16782;
	#10 counter$count = 16783;
	#10 counter$count = 16784;
	#10 counter$count = 16785;
	#10 counter$count = 16786;
	#10 counter$count = 16787;
	#10 counter$count = 16788;
	#10 counter$count = 16789;
	#10 counter$count = 16790;
	#10 counter$count = 16791;
	#10 counter$count = 16792;
	#10 counter$count = 16793;
	#10 counter$count = 16794;
	#10 counter$count = 16795;
	#10 counter$count = 16796;
	#10 counter$count = 16797;
	#10 counter$count = 16798;
	#10 counter$count = 16799;
	#10 counter$count = 16800;
	#10 counter$count = 16801;
	#10 counter$count = 16802;
	#10 counter$count = 16803;
	#10 counter$count = 16804;
	#10 counter$count = 16805;
	#10 counter$count = 16806;
	#10 counter$count = 16807;
	#10 counter$count = 16808;
	#10 counter$count = 16809;
	#10 counter$count = 16810;
	#10 counter$count = 16811;
	#10 counter$count = 16812;
	#10 counter$count = 16813;
	#10 counter$count = 16814;
	#10 counter$count = 16815;
	#10 counter$count = 16816;
	#10 counter$count = 16817;
	#10 counter$count = 16818;
	#10 counter$count = 16819;
	#10 counter$count = 16820;
	#10 counter$count = 16821;
	#10 counter$count = 16822;
	#10 counter$count = 16823;
	#10 counter$count = 16824;
	#10 counter$count = 16825;
	#10 counter$count = 16826;
	#10 counter$count = 16827;
	#10 counter$count = 16828;
	#10 counter$count = 16829;
	#10 counter$count = 16830;
	#10 counter$count = 16831;
	#10 counter$count = 16832;
	#10 counter$count = 16833;
	#10 counter$count = 16834;
	#10 counter$count = 16835;
	#10 counter$count = 16836;
	#10 counter$count = 16837;
	#10 counter$count = 16838;
	#10 counter$count = 16839;
	#10 counter$count = 16840;
	#10 counter$count = 16841;
	#10 counter$count = 16842;
	#10 counter$count = 16843;
	#10 counter$count = 16844;
	#10 counter$count = 16845;
	#10 counter$count = 16846;
	#10 counter$count = 16847;
	#10 counter$count = 16848;
	#10 counter$count = 16849;
	#10 counter$count = 16850;
	#10 counter$count = 16851;
	#10 counter$count = 16852;
	#10 counter$count = 16853;
	#10 counter$count = 16854;
	#10 counter$count = 16855;
	#10 counter$count = 16856;
	#10 counter$count = 16857;
	#10 counter$count = 16858;
	#10 counter$count = 16859;
	#10 counter$count = 16860;
	#10 counter$count = 16861;
	#10 counter$count = 16862;
	#10 counter$count = 16863;
	#10 counter$count = 16864;
	#10 counter$count = 16865;
	#10 counter$count = 16866;
	#10 counter$count = 16867;
	#10 counter$count = 16868;
	#10 counter$count = 16869;
	#10 counter$count = 16870;
	#10 counter$count = 16871;
	#10 counter$count = 16872;
	#10 counter$count = 16873;
	#10 counter$count = 16874;
	#10 counter$count = 16875;
	#10 counter$count = 16876;
	#10 counter$count = 16877;
	#10 counter$count = 16878;
	#10 counter$count = 16879;
	#10 counter$count = 16880;
	#10 counter$count = 16881;
	#10 counter$count = 16882;
	#10 counter$count = 16883;
	#10 counter$count = 16884;
	#10 counter$count = 16885;
	#10 counter$count = 16886;
	#10 counter$count = 16887;
	#10 counter$count = 16888;
	#10 counter$count = 16889;
	#10 counter$count = 16890;
	#10 counter$count = 16891;
	#10 counter$count = 16892;
	#10 counter$count = 16893;
	#10 counter$count = 16894;
	#10 counter$count = 16895;
	#10 counter$count = 16896;
	#10 counter$count = 16897;
	#10 counter$count = 16898;
	#10 counter$count = 16899;
	#10 counter$count = 16900;
	#10 counter$count = 16901;
	#10 counter$count = 16902;
	#10 counter$count = 16903;
	#10 counter$count = 16904;
	#10 counter$count = 16905;
	#10 counter$count = 16906;
	#10 counter$count = 16907;
	#10 counter$count = 16908;
	#10 counter$count = 16909;
	#10 counter$count = 16910;
	#10 counter$count = 16911;
	#10 counter$count = 16912;
	#10 counter$count = 16913;
	#10 counter$count = 16914;
	#10 counter$count = 16915;
	#10 counter$count = 16916;
	#10 counter$count = 16917;
	#10 counter$count = 16918;
	#10 counter$count = 16919;
	#10 counter$count = 16920;
	#10 counter$count = 16921;
	#10 counter$count = 16922;
	#10 counter$count = 16923;
	#10 counter$count = 16924;
	#10 counter$count = 16925;
	#10 counter$count = 16926;
	#10 counter$count = 16927;
	#10 counter$count = 16928;
	#10 counter$count = 16929;
	#10 counter$count = 16930;
	#10 counter$count = 16931;
	#10 counter$count = 16932;
	#10 counter$count = 16933;
	#10 counter$count = 16934;
	#10 counter$count = 16935;
	#10 counter$count = 16936;
	#10 counter$count = 16937;
	#10 counter$count = 16938;
	#10 counter$count = 16939;
	#10 counter$count = 16940;
	#10 counter$count = 16941;
	#10 counter$count = 16942;
	#10 counter$count = 16943;
	#10 counter$count = 16944;
	#10 counter$count = 16945;
	#10 counter$count = 16946;
	#10 counter$count = 16947;
	#10 counter$count = 16948;
	#10 counter$count = 16949;
	#10 counter$count = 16950;
	#10 counter$count = 16951;
	#10 counter$count = 16952;
	#10 counter$count = 16953;
	#10 counter$count = 16954;
	#10 counter$count = 16955;
	#10 counter$count = 16956;
	#10 counter$count = 16957;
	#10 counter$count = 16958;
	#10 counter$count = 16959;
	#10 counter$count = 16960;
	#10 counter$count = 16961;
	#10 counter$count = 16962;
	#10 counter$count = 16963;
	#10 counter$count = 16964;
	#10 counter$count = 16965;
	#10 counter$count = 16966;
	#10 counter$count = 16967;
	#10 counter$count = 16968;
	#10 counter$count = 16969;
	#10 counter$count = 16970;
	#10 counter$count = 16971;
	#10 counter$count = 16972;
	#10 counter$count = 16973;
	#10 counter$count = 16974;
	#10 counter$count = 16975;
	#10 counter$count = 16976;
	#10 counter$count = 16977;
	#10 counter$count = 16978;
	#10 counter$count = 16979;
	#10 counter$count = 16980;
	#10 counter$count = 16981;
	#10 counter$count = 16982;
	#10 counter$count = 16983;
	#10 counter$count = 16984;
	#10 counter$count = 16985;
	#10 counter$count = 16986;
	#10 counter$count = 16987;
	#10 counter$count = 16988;
	#10 counter$count = 16989;
	#10 counter$count = 16990;
	#10 counter$count = 16991;
	#10 counter$count = 16992;
	#10 counter$count = 16993;
	#10 counter$count = 16994;
	#10 counter$count = 16995;
	#10 counter$count = 16996;
	#10 counter$count = 16997;
	#10 counter$count = 16998;
	#10 counter$count = 16999;
	#10 counter$count = 17000;
	#10 counter$count = 17001;
	#10 counter$count = 17002;
	#10 counter$count = 17003;
	#10 counter$count = 17004;
	#10 counter$count = 17005;
	#10 counter$count = 17006;
	#10 counter$count = 17007;
	#10 counter$count = 17008;
	#10 counter$count = 17009;
	#10 counter$count = 17010;
	#10 counter$count = 17011;
	#10 counter$count = 17012;
	#10 counter$count = 17013;
	#10 counter$count = 17014;
	#10 counter$count = 17015;
	#10 counter$count = 17016;
	#10 counter$count = 17017;
	#10 counter$count = 17018;
	#10 counter$count = 17019;
	#10 counter$count = 17020;
	#10 counter$count = 17021;
	#10 counter$count = 17022;
	#10 counter$count = 17023;
	#10 counter$count = 17024;
	#10 counter$count = 17025;
	#10 counter$count = 17026;
	#10 counter$count = 17027;
	#10 counter$count = 17028;
	#10 counter$count = 17029;
	#10 counter$count = 17030;
	#10 counter$count = 17031;
	#10 counter$count = 17032;
	#10 counter$count = 17033;
	#10 counter$count = 17034;
	#10 counter$count = 17035;
	#10 counter$count = 17036;
	#10 counter$count = 17037;
	#10 counter$count = 17038;
	#10 counter$count = 17039;
	#10 counter$count = 17040;
	#10 counter$count = 17041;
	#10 counter$count = 17042;
	#10 counter$count = 17043;
	#10 counter$count = 17044;
	#10 counter$count = 17045;
	#10 counter$count = 17046;
	#10 counter$count = 17047;
	#10 counter$count = 17048;
	#10 counter$count = 17049;
	#10 counter$count = 17050;
	#10 counter$count = 17051;
	#10 counter$count = 17052;
	#10 counter$count = 17053;
	#10 counter$count = 17054;
	#10 counter$count = 17055;
	#10 counter$count = 17056;
	#10 counter$count = 17057;
	#10 counter$count = 17058;
	#10 counter$count = 17059;
	#10 counter$count = 17060;
	#10 counter$count = 17061;
	#10 counter$count = 17062;
	#10 counter$count = 17063;
	#10 counter$count = 17064;
	#10 counter$count = 17065;
	#10 counter$count = 17066;
	#10 counter$count = 17067;
	#10 counter$count = 17068;
	#10 counter$count = 17069;
	#10 counter$count = 17070;
	#10 counter$count = 17071;
	#10 counter$count = 17072;
	#10 counter$count = 17073;
	#10 counter$count = 17074;
	#10 counter$count = 17075;
	#10 counter$count = 17076;
	#10 counter$count = 17077;
	#10 counter$count = 17078;
	#10 counter$count = 17079;
	#10 counter$count = 17080;
	#10 counter$count = 17081;
	#10 counter$count = 17082;
	#10 counter$count = 17083;
	#10 counter$count = 17084;
	#10 counter$count = 17085;
	#10 counter$count = 17086;
	#10 counter$count = 17087;
	#10 counter$count = 17088;
	#10 counter$count = 17089;
	#10 counter$count = 17090;
	#10 counter$count = 17091;
	#10 counter$count = 17092;
	#10 counter$count = 17093;
	#10 counter$count = 17094;
	#10 counter$count = 17095;
	#10 counter$count = 17096;
	#10 counter$count = 17097;
	#10 counter$count = 17098;
	#10 counter$count = 17099;
	#10 counter$count = 17100;
	#10 counter$count = 17101;
	#10 counter$count = 17102;
	#10 counter$count = 17103;
	#10 counter$count = 17104;
	#10 counter$count = 17105;
	#10 counter$count = 17106;
	#10 counter$count = 17107;
	#10 counter$count = 17108;
	#10 counter$count = 17109;
	#10 counter$count = 17110;
	#10 counter$count = 17111;
	#10 counter$count = 17112;
	#10 counter$count = 17113;
	#10 counter$count = 17114;
	#10 counter$count = 17115;
	#10 counter$count = 17116;
	#10 counter$count = 17117;
	#10 counter$count = 17118;
	#10 counter$count = 17119;
	#10 counter$count = 17120;
	#10 counter$count = 17121;
	#10 counter$count = 17122;
	#10 counter$count = 17123;
	#10 counter$count = 17124;
	#10 counter$count = 17125;
	#10 counter$count = 17126;
	#10 counter$count = 17127;
	#10 counter$count = 17128;
	#10 counter$count = 17129;
	#10 counter$count = 17130;
	#10 counter$count = 17131;
	#10 counter$count = 17132;
	#10 counter$count = 17133;
	#10 counter$count = 17134;
	#10 counter$count = 17135;
	#10 counter$count = 17136;
	#10 counter$count = 17137;
	#10 counter$count = 17138;
	#10 counter$count = 17139;
	#10 counter$count = 17140;
	#10 counter$count = 17141;
	#10 counter$count = 17142;
	#10 counter$count = 17143;
	#10 counter$count = 17144;
	#10 counter$count = 17145;
	#10 counter$count = 17146;
	#10 counter$count = 17147;
	#10 counter$count = 17148;
	#10 counter$count = 17149;
	#10 counter$count = 17150;
	#10 counter$count = 17151;
	#10 counter$count = 17152;
	#10 counter$count = 17153;
	#10 counter$count = 17154;
	#10 counter$count = 17155;
	#10 counter$count = 17156;
	#10 counter$count = 17157;
	#10 counter$count = 17158;
	#10 counter$count = 17159;
	#10 counter$count = 17160;
	#10 counter$count = 17161;
	#10 counter$count = 17162;
	#10 counter$count = 17163;
	#10 counter$count = 17164;
	#10 counter$count = 17165;
	#10 counter$count = 17166;
	#10 counter$count = 17167;
	#10 counter$count = 17168;
	#10 counter$count = 17169;
	#10 counter$count = 17170;
	#10 counter$count = 17171;
	#10 counter$count = 17172;
	#10 counter$count = 17173;
	#10 counter$count = 17174;
	#10 counter$count = 17175;
	#10 counter$count = 17176;
	#10 counter$count = 17177;
	#10 counter$count = 17178;
	#10 counter$count = 17179;
	#10 counter$count = 17180;
	#10 counter$count = 17181;
	#10 counter$count = 17182;
	#10 counter$count = 17183;
	#10 counter$count = 17184;
	#10 counter$count = 17185;
	#10 counter$count = 17186;
	#10 counter$count = 17187;
	#10 counter$count = 17188;
	#10 counter$count = 17189;
	#10 counter$count = 17190;
	#10 counter$count = 17191;
	#10 counter$count = 17192;
	#10 counter$count = 17193;
	#10 counter$count = 17194;
	#10 counter$count = 17195;
	#10 counter$count = 17196;
	#10 counter$count = 17197;
	#10 counter$count = 17198;
	#10 counter$count = 17199;
	#10 counter$count = 17200;
	#10 counter$count = 17201;
	#10 counter$count = 17202;
	#10 counter$count = 17203;
	#10 counter$count = 17204;
	#10 counter$count = 17205;
	#10 counter$count = 17206;
	#10 counter$count = 17207;
	#10 counter$count = 17208;
	#10 counter$count = 17209;
	#10 counter$count = 17210;
	#10 counter$count = 17211;
	#10 counter$count = 17212;
	#10 counter$count = 17213;
	#10 counter$count = 17214;
	#10 counter$count = 17215;
	#10 counter$count = 17216;
	#10 counter$count = 17217;
	#10 counter$count = 17218;
	#10 counter$count = 17219;
	#10 counter$count = 17220;
	#10 counter$count = 17221;
	#10 counter$count = 17222;
	#10 counter$count = 17223;
	#10 counter$count = 17224;
	#10 counter$count = 17225;
	#10 counter$count = 17226;
	#10 counter$count = 17227;
	#10 counter$count = 17228;
	#10 counter$count = 17229;
	#10 counter$count = 17230;
	#10 counter$count = 17231;
	#10 counter$count = 17232;
	#10 counter$count = 17233;
	#10 counter$count = 17234;
	#10 counter$count = 17235;
	#10 counter$count = 17236;
	#10 counter$count = 17237;
	#10 counter$count = 17238;
	#10 counter$count = 17239;
	#10 counter$count = 17240;
	#10 counter$count = 17241;
	#10 counter$count = 17242;
	#10 counter$count = 17243;
	#10 counter$count = 17244;
	#10 counter$count = 17245;
	#10 counter$count = 17246;
	#10 counter$count = 17247;
	#10 counter$count = 17248;
	#10 counter$count = 17249;
	#10 counter$count = 17250;
	#10 counter$count = 17251;
	#10 counter$count = 17252;
	#10 counter$count = 17253;
	#10 counter$count = 17254;
	#10 counter$count = 17255;
	#10 counter$count = 17256;
	#10 counter$count = 17257;
	#10 counter$count = 17258;
	#10 counter$count = 17259;
	#10 counter$count = 17260;
	#10 counter$count = 17261;
	#10 counter$count = 17262;
	#10 counter$count = 17263;
	#10 counter$count = 17264;
	#10 counter$count = 17265;
	#10 counter$count = 17266;
	#10 counter$count = 17267;
	#10 counter$count = 17268;
	#10 counter$count = 17269;
	#10 counter$count = 17270;
	#10 counter$count = 17271;
	#10 counter$count = 17272;
	#10 counter$count = 17273;
	#10 counter$count = 17274;
	#10 counter$count = 17275;
	#10 counter$count = 17276;
	#10 counter$count = 17277;
	#10 counter$count = 17278;
	#10 counter$count = 17279;
	#10 counter$count = 17280;
	#10 counter$count = 17281;
	#10 counter$count = 17282;
	#10 counter$count = 17283;
	#10 counter$count = 17284;
	#10 counter$count = 17285;
	#10 counter$count = 17286;
	#10 counter$count = 17287;
	#10 counter$count = 17288;
	#10 counter$count = 17289;
	#10 counter$count = 17290;
	#10 counter$count = 17291;
	#10 counter$count = 17292;
	#10 counter$count = 17293;
	#10 counter$count = 17294;
	#10 counter$count = 17295;
	#10 counter$count = 17296;
	#10 counter$count = 17297;
	#10 counter$count = 17298;
	#10 counter$count = 17299;
	#10 counter$count = 17300;
	#10 counter$count = 17301;
	#10 counter$count = 17302;
	#10 counter$count = 17303;
	#10 counter$count = 17304;
	#10 counter$count = 17305;
	#10 counter$count = 17306;
	#10 counter$count = 17307;
	#10 counter$count = 17308;
	#10 counter$count = 17309;
	#10 counter$count = 17310;
	#10 counter$count = 17311;
	#10 counter$count = 17312;
	#10 counter$count = 17313;
	#10 counter$count = 17314;
	#10 counter$count = 17315;
	#10 counter$count = 17316;
	#10 counter$count = 17317;
	#10 counter$count = 17318;
	#10 counter$count = 17319;
	#10 counter$count = 17320;
	#10 counter$count = 17321;
	#10 counter$count = 17322;
	#10 counter$count = 17323;
	#10 counter$count = 17324;
	#10 counter$count = 17325;
	#10 counter$count = 17326;
	#10 counter$count = 17327;
	#10 counter$count = 17328;
	#10 counter$count = 17329;
	#10 counter$count = 17330;
	#10 counter$count = 17331;
	#10 counter$count = 17332;
	#10 counter$count = 17333;
	#10 counter$count = 17334;
	#10 counter$count = 17335;
	#10 counter$count = 17336;
	#10 counter$count = 17337;
	#10 counter$count = 17338;
	#10 counter$count = 17339;
	#10 counter$count = 17340;
	#10 counter$count = 17341;
	#10 counter$count = 17342;
	#10 counter$count = 17343;
	#10 counter$count = 17344;
	#10 counter$count = 17345;
	#10 counter$count = 17346;
	#10 counter$count = 17347;
	#10 counter$count = 17348;
	#10 counter$count = 17349;
	#10 counter$count = 17350;
	#10 counter$count = 17351;
	#10 counter$count = 17352;
	#10 counter$count = 17353;
	#10 counter$count = 17354;
	#10 counter$count = 17355;
	#10 counter$count = 17356;
	#10 counter$count = 17357;
	#10 counter$count = 17358;
	#10 counter$count = 17359;
	#10 counter$count = 17360;
	#10 counter$count = 17361;
	#10 counter$count = 17362;
	#10 counter$count = 17363;
	#10 counter$count = 17364;
	#10 counter$count = 17365;
	#10 counter$count = 17366;
	#10 counter$count = 17367;
	#10 counter$count = 17368;
	#10 counter$count = 17369;
	#10 counter$count = 17370;
	#10 counter$count = 17371;
	#10 counter$count = 17372;
	#10 counter$count = 17373;
	#10 counter$count = 17374;
	#10 counter$count = 17375;
	#10 counter$count = 17376;
	#10 counter$count = 17377;
	#10 counter$count = 17378;
	#10 counter$count = 17379;
	#10 counter$count = 17380;
	#10 counter$count = 17381;
	#10 counter$count = 17382;
	#10 counter$count = 17383;
	#10 counter$count = 17384;
	#10 counter$count = 17385;
	#10 counter$count = 17386;
	#10 counter$count = 17387;
	#10 counter$count = 17388;
	#10 counter$count = 17389;
	#10 counter$count = 17390;
	#10 counter$count = 17391;
	#10 counter$count = 17392;
	#10 counter$count = 17393;
	#10 counter$count = 17394;
	#10 counter$count = 17395;
	#10 counter$count = 17396;
	#10 counter$count = 17397;
	#10 counter$count = 17398;
	#10 counter$count = 17399;
	#10 counter$count = 17400;
	#10 counter$count = 17401;
	#10 counter$count = 17402;
	#10 counter$count = 17403;
	#10 counter$count = 17404;
	#10 counter$count = 17405;
	#10 counter$count = 17406;
	#10 counter$count = 17407;
	#10 counter$count = 17408;
	#10 counter$count = 17409;
	#10 counter$count = 17410;
	#10 counter$count = 17411;
	#10 counter$count = 17412;
	#10 counter$count = 17413;
	#10 counter$count = 17414;
	#10 counter$count = 17415;
	#10 counter$count = 17416;
	#10 counter$count = 17417;
	#10 counter$count = 17418;
	#10 counter$count = 17419;
	#10 counter$count = 17420;
	#10 counter$count = 17421;
	#10 counter$count = 17422;
	#10 counter$count = 17423;
	#10 counter$count = 17424;
	#10 counter$count = 17425;
	#10 counter$count = 17426;
	#10 counter$count = 17427;
	#10 counter$count = 17428;
	#10 counter$count = 17429;
	#10 counter$count = 17430;
	#10 counter$count = 17431;
	#10 counter$count = 17432;
	#10 counter$count = 17433;
	#10 counter$count = 17434;
	#10 counter$count = 17435;
	#10 counter$count = 17436;
	#10 counter$count = 17437;
	#10 counter$count = 17438;
	#10 counter$count = 17439;
	#10 counter$count = 17440;
	#10 counter$count = 17441;
	#10 counter$count = 17442;
	#10 counter$count = 17443;
	#10 counter$count = 17444;
	#10 counter$count = 17445;
	#10 counter$count = 17446;
	#10 counter$count = 17447;
	#10 counter$count = 17448;
	#10 counter$count = 17449;
	#10 counter$count = 17450;
	#10 counter$count = 17451;
	#10 counter$count = 17452;
	#10 counter$count = 17453;
	#10 counter$count = 17454;
	#10 counter$count = 17455;
	#10 counter$count = 17456;
	#10 counter$count = 17457;
	#10 counter$count = 17458;
	#10 counter$count = 17459;
	#10 counter$count = 17460;
	#10 counter$count = 17461;
	#10 counter$count = 17462;
	#10 counter$count = 17463;
	#10 counter$count = 17464;
	#10 counter$count = 17465;
	#10 counter$count = 17466;
	#10 counter$count = 17467;
	#10 counter$count = 17468;
	#10 counter$count = 17469;
	#10 counter$count = 17470;
	#10 counter$count = 17471;
	#10 counter$count = 17472;
	#10 counter$count = 17473;
	#10 counter$count = 17474;
	#10 counter$count = 17475;
	#10 counter$count = 17476;
	#10 counter$count = 17477;
	#10 counter$count = 17478;
	#10 counter$count = 17479;
	#10 counter$count = 17480;
	#10 counter$count = 17481;
	#10 counter$count = 17482;
	#10 counter$count = 17483;
	#10 counter$count = 17484;
	#10 counter$count = 17485;
	#10 counter$count = 17486;
	#10 counter$count = 17487;
	#10 counter$count = 17488;
	#10 counter$count = 17489;
	#10 counter$count = 17490;
	#10 counter$count = 17491;
	#10 counter$count = 17492;
	#10 counter$count = 17493;
	#10 counter$count = 17494;
	#10 counter$count = 17495;
	#10 counter$count = 17496;
	#10 counter$count = 17497;
	#10 counter$count = 17498;
	#10 counter$count = 17499;
	#10 counter$count = 17500;
	#10 counter$count = 17501;
	#10 counter$count = 17502;
	#10 counter$count = 17503;
	#10 counter$count = 17504;
	#10 counter$count = 17505;
	#10 counter$count = 17506;
	#10 counter$count = 17507;
	#10 counter$count = 17508;
	#10 counter$count = 17509;
	#10 counter$count = 17510;
	#10 counter$count = 17511;
	#10 counter$count = 17512;
	#10 counter$count = 17513;
	#10 counter$count = 17514;
	#10 counter$count = 17515;
	#10 counter$count = 17516;
	#10 counter$count = 17517;
	#10 counter$count = 17518;
	#10 counter$count = 17519;
	#10 counter$count = 17520;
	#10 counter$count = 17521;
	#10 counter$count = 17522;
	#10 counter$count = 17523;
	#10 counter$count = 17524;
	#10 counter$count = 17525;
	#10 counter$count = 17526;
	#10 counter$count = 17527;
	#10 counter$count = 17528;
	#10 counter$count = 17529;
	#10 counter$count = 17530;
	#10 counter$count = 17531;
	#10 counter$count = 17532;
	#10 counter$count = 17533;
	#10 counter$count = 17534;
	#10 counter$count = 17535;
	#10 counter$count = 17536;
	#10 counter$count = 17537;
	#10 counter$count = 17538;
	#10 counter$count = 17539;
	#10 counter$count = 17540;
	#10 counter$count = 17541;
	#10 counter$count = 17542;
	#10 counter$count = 17543;
	#10 counter$count = 17544;
	#10 counter$count = 17545;
	#10 counter$count = 17546;
	#10 counter$count = 17547;
	#10 counter$count = 17548;
	#10 counter$count = 17549;
	#10 counter$count = 17550;
	#10 counter$count = 17551;
	#10 counter$count = 17552;
	#10 counter$count = 17553;
	#10 counter$count = 17554;
	#10 counter$count = 17555;
	#10 counter$count = 17556;
	#10 counter$count = 17557;
	#10 counter$count = 17558;
	#10 counter$count = 17559;
	#10 counter$count = 17560;
	#10 counter$count = 17561;
	#10 counter$count = 17562;
	#10 counter$count = 17563;
	#10 counter$count = 17564;
	#10 counter$count = 17565;
	#10 counter$count = 17566;
	#10 counter$count = 17567;
	#10 counter$count = 17568;
	#10 counter$count = 17569;
	#10 counter$count = 17570;
	#10 counter$count = 17571;
	#10 counter$count = 17572;
	#10 counter$count = 17573;
	#10 counter$count = 17574;
	#10 counter$count = 17575;
	#10 counter$count = 17576;
	#10 counter$count = 17577;
	#10 counter$count = 17578;
	#10 counter$count = 17579;
	#10 counter$count = 17580;
	#10 counter$count = 17581;
	#10 counter$count = 17582;
	#10 counter$count = 17583;
	#10 counter$count = 17584;
	#10 counter$count = 17585;
	#10 counter$count = 17586;
	#10 counter$count = 17587;
	#10 counter$count = 17588;
	#10 counter$count = 17589;
	#10 counter$count = 17590;
	#10 counter$count = 17591;
	#10 counter$count = 17592;
	#10 counter$count = 17593;
	#10 counter$count = 17594;
	#10 counter$count = 17595;
	#10 counter$count = 17596;
	#10 counter$count = 17597;
	#10 counter$count = 17598;
	#10 counter$count = 17599;
	#10 counter$count = 17600;
	#10 counter$count = 17601;
	#10 counter$count = 17602;
	#10 counter$count = 17603;
	#10 counter$count = 17604;
	#10 counter$count = 17605;
	#10 counter$count = 17606;
	#10 counter$count = 17607;
	#10 counter$count = 17608;
	#10 counter$count = 17609;
	#10 counter$count = 17610;
	#10 counter$count = 17611;
	#10 counter$count = 17612;
	#10 counter$count = 17613;
	#10 counter$count = 17614;
	#10 counter$count = 17615;
	#10 counter$count = 17616;
	#10 counter$count = 17617;
	#10 counter$count = 17618;
	#10 counter$count = 17619;
	#10 counter$count = 17620;
	#10 counter$count = 17621;
	#10 counter$count = 17622;
	#10 counter$count = 17623;
	#10 counter$count = 17624;
	#10 counter$count = 17625;
	#10 counter$count = 17626;
	#10 counter$count = 17627;
	#10 counter$count = 17628;
	#10 counter$count = 17629;
	#10 counter$count = 17630;
	#10 counter$count = 17631;
	#10 counter$count = 17632;
	#10 counter$count = 17633;
	#10 counter$count = 17634;
	#10 counter$count = 17635;
	#10 counter$count = 17636;
	#10 counter$count = 17637;
	#10 counter$count = 17638;
	#10 counter$count = 17639;
	#10 counter$count = 17640;
	#10 counter$count = 17641;
	#10 counter$count = 17642;
	#10 counter$count = 17643;
	#10 counter$count = 17644;
	#10 counter$count = 17645;
	#10 counter$count = 17646;
	#10 counter$count = 17647;
	#10 counter$count = 17648;
	#10 counter$count = 17649;
	#10 counter$count = 17650;
	#10 counter$count = 17651;
	#10 counter$count = 17652;
	#10 counter$count = 17653;
	#10 counter$count = 17654;
	#10 counter$count = 17655;
	#10 counter$count = 17656;
	#10 counter$count = 17657;
	#10 counter$count = 17658;
	#10 counter$count = 17659;
	#10 counter$count = 17660;
	#10 counter$count = 17661;
	#10 counter$count = 17662;
	#10 counter$count = 17663;
	#10 counter$count = 17664;
	#10 counter$count = 17665;
	#10 counter$count = 17666;
	#10 counter$count = 17667;
	#10 counter$count = 17668;
	#10 counter$count = 17669;
	#10 counter$count = 17670;
	#10 counter$count = 17671;
	#10 counter$count = 17672;
	#10 counter$count = 17673;
	#10 counter$count = 17674;
	#10 counter$count = 17675;
	#10 counter$count = 17676;
	#10 counter$count = 17677;
	#10 counter$count = 17678;
	#10 counter$count = 17679;
	#10 counter$count = 17680;
	#10 counter$count = 17681;
	#10 counter$count = 17682;
	#10 counter$count = 17683;
	#10 counter$count = 17684;
	#10 counter$count = 17685;
	#10 counter$count = 17686;
	#10 counter$count = 17687;
	#10 counter$count = 17688;
	#10 counter$count = 17689;
	#10 counter$count = 17690;
	#10 counter$count = 17691;
	#10 counter$count = 17692;
	#10 counter$count = 17693;
	#10 counter$count = 17694;
	#10 counter$count = 17695;
	#10 counter$count = 17696;
	#10 counter$count = 17697;
	#10 counter$count = 17698;
	#10 counter$count = 17699;
	#10 counter$count = 17700;
	#10 counter$count = 17701;
	#10 counter$count = 17702;
	#10 counter$count = 17703;
	#10 counter$count = 17704;
	#10 counter$count = 17705;
	#10 counter$count = 17706;
	#10 counter$count = 17707;
	#10 counter$count = 17708;
	#10 counter$count = 17709;
	#10 counter$count = 17710;
	#10 counter$count = 17711;
	#10 counter$count = 17712;
	#10 counter$count = 17713;
	#10 counter$count = 17714;
	#10 counter$count = 17715;
	#10 counter$count = 17716;
	#10 counter$count = 17717;
	#10 counter$count = 17718;
	#10 counter$count = 17719;
	#10 counter$count = 17720;
	#10 counter$count = 17721;
	#10 counter$count = 17722;
	#10 counter$count = 17723;
	#10 counter$count = 17724;
	#10 counter$count = 17725;
	#10 counter$count = 17726;
	#10 counter$count = 17727;
	#10 counter$count = 17728;
	#10 counter$count = 17729;
	#10 counter$count = 17730;
	#10 counter$count = 17731;
	#10 counter$count = 17732;
	#10 counter$count = 17733;
	#10 counter$count = 17734;
	#10 counter$count = 17735;
	#10 counter$count = 17736;
	#10 counter$count = 17737;
	#10 counter$count = 17738;
	#10 counter$count = 17739;
	#10 counter$count = 17740;
	#10 counter$count = 17741;
	#10 counter$count = 17742;
	#10 counter$count = 17743;
	#10 counter$count = 17744;
	#10 counter$count = 17745;
	#10 counter$count = 17746;
	#10 counter$count = 17747;
	#10 counter$count = 17748;
	#10 counter$count = 17749;
	#10 counter$count = 17750;
	#10 counter$count = 17751;
	#10 counter$count = 17752;
	#10 counter$count = 17753;
	#10 counter$count = 17754;
	#10 counter$count = 17755;
	#10 counter$count = 17756;
	#10 counter$count = 17757;
	#10 counter$count = 17758;
	#10 counter$count = 17759;
	#10 counter$count = 17760;
	#10 counter$count = 17761;
	#10 counter$count = 17762;
	#10 counter$count = 17763;
	#10 counter$count = 17764;
	#10 counter$count = 17765;
	#10 counter$count = 17766;
	#10 counter$count = 17767;
	#10 counter$count = 17768;
	#10 counter$count = 17769;
	#10 counter$count = 17770;
	#10 counter$count = 17771;
	#10 counter$count = 17772;
	#10 counter$count = 17773;
	#10 counter$count = 17774;
	#10 counter$count = 17775;
	#10 counter$count = 17776;
	#10 counter$count = 17777;
	#10 counter$count = 17778;
	#10 counter$count = 17779;
	#10 counter$count = 17780;
	#10 counter$count = 17781;
	#10 counter$count = 17782;
	#10 counter$count = 17783;
	#10 counter$count = 17784;
	#10 counter$count = 17785;
	#10 counter$count = 17786;
	#10 counter$count = 17787;
	#10 counter$count = 17788;
	#10 counter$count = 17789;
	#10 counter$count = 17790;
	#10 counter$count = 17791;
	#10 counter$count = 17792;
	#10 counter$count = 17793;
	#10 counter$count = 17794;
	#10 counter$count = 17795;
	#10 counter$count = 17796;
	#10 counter$count = 17797;
	#10 counter$count = 17798;
	#10 counter$count = 17799;
	#10 counter$count = 17800;
	#10 counter$count = 17801;
	#10 counter$count = 17802;
	#10 counter$count = 17803;
	#10 counter$count = 17804;
	#10 counter$count = 17805;
	#10 counter$count = 17806;
	#10 counter$count = 17807;
	#10 counter$count = 17808;
	#10 counter$count = 17809;
	#10 counter$count = 17810;
	#10 counter$count = 17811;
	#10 counter$count = 17812;
	#10 counter$count = 17813;
	#10 counter$count = 17814;
	#10 counter$count = 17815;
	#10 counter$count = 17816;
	#10 counter$count = 17817;
	#10 counter$count = 17818;
	#10 counter$count = 17819;
	#10 counter$count = 17820;
	#10 counter$count = 17821;
	#10 counter$count = 17822;
	#10 counter$count = 17823;
	#10 counter$count = 17824;
	#10 counter$count = 17825;
	#10 counter$count = 17826;
	#10 counter$count = 17827;
	#10 counter$count = 17828;
	#10 counter$count = 17829;
	#10 counter$count = 17830;
	#10 counter$count = 17831;
	#10 counter$count = 17832;
	#10 counter$count = 17833;
	#10 counter$count = 17834;
	#10 counter$count = 17835;
	#10 counter$count = 17836;
	#10 counter$count = 17837;
	#10 counter$count = 17838;
	#10 counter$count = 17839;
	#10 counter$count = 17840;
	#10 counter$count = 17841;
	#10 counter$count = 17842;
	#10 counter$count = 17843;
	#10 counter$count = 17844;
	#10 counter$count = 17845;
	#10 counter$count = 17846;
	#10 counter$count = 17847;
	#10 counter$count = 17848;
	#10 counter$count = 17849;
	#10 counter$count = 17850;
	#10 counter$count = 17851;
	#10 counter$count = 17852;
	#10 counter$count = 17853;
	#10 counter$count = 17854;
	#10 counter$count = 17855;
	#10 counter$count = 17856;
	#10 counter$count = 17857;
	#10 counter$count = 17858;
	#10 counter$count = 17859;
	#10 counter$count = 17860;
	#10 counter$count = 17861;
	#10 counter$count = 17862;
	#10 counter$count = 17863;
	#10 counter$count = 17864;
	#10 counter$count = 17865;
	#10 counter$count = 17866;
	#10 counter$count = 17867;
	#10 counter$count = 17868;
	#10 counter$count = 17869;
	#10 counter$count = 17870;
	#10 counter$count = 17871;
	#10 counter$count = 17872;
	#10 counter$count = 17873;
	#10 counter$count = 17874;
	#10 counter$count = 17875;
	#10 counter$count = 17876;
	#10 counter$count = 17877;
	#10 counter$count = 17878;
	#10 counter$count = 17879;
	#10 counter$count = 17880;
	#10 counter$count = 17881;
	#10 counter$count = 17882;
	#10 counter$count = 17883;
	#10 counter$count = 17884;
	#10 counter$count = 17885;
	#10 counter$count = 17886;
	#10 counter$count = 17887;
	#10 counter$count = 17888;
	#10 counter$count = 17889;
	#10 counter$count = 17890;
	#10 counter$count = 17891;
	#10 counter$count = 17892;
	#10 counter$count = 17893;
	#10 counter$count = 17894;
	#10 counter$count = 17895;
	#10 counter$count = 17896;
	#10 counter$count = 17897;
	#10 counter$count = 17898;
	#10 counter$count = 17899;
	#10 counter$count = 17900;
	#10 counter$count = 17901;
	#10 counter$count = 17902;
	#10 counter$count = 17903;
	#10 counter$count = 17904;
	#10 counter$count = 17905;
	#10 counter$count = 17906;
	#10 counter$count = 17907;
	#10 counter$count = 17908;
	#10 counter$count = 17909;
	#10 counter$count = 17910;
	#10 counter$count = 17911;
	#10 counter$count = 17912;
	#10 counter$count = 17913;
	#10 counter$count = 17914;
	#10 counter$count = 17915;
	#10 counter$count = 17916;
	#10 counter$count = 17917;
	#10 counter$count = 17918;
	#10 counter$count = 17919;
	#10 counter$count = 17920;
	#10 counter$count = 17921;
	#10 counter$count = 17922;
	#10 counter$count = 17923;
	#10 counter$count = 17924;
	#10 counter$count = 17925;
	#10 counter$count = 17926;
	#10 counter$count = 17927;
	#10 counter$count = 17928;
	#10 counter$count = 17929;
	#10 counter$count = 17930;
	#10 counter$count = 17931;
	#10 counter$count = 17932;
	#10 counter$count = 17933;
	#10 counter$count = 17934;
	#10 counter$count = 17935;
	#10 counter$count = 17936;
	#10 counter$count = 17937;
	#10 counter$count = 17938;
	#10 counter$count = 17939;
	#10 counter$count = 17940;
	#10 counter$count = 17941;
	#10 counter$count = 17942;
	#10 counter$count = 17943;
	#10 counter$count = 17944;
	#10 counter$count = 17945;
	#10 counter$count = 17946;
	#10 counter$count = 17947;
	#10 counter$count = 17948;
	#10 counter$count = 17949;
	#10 counter$count = 17950;
	#10 counter$count = 17951;
	#10 counter$count = 17952;
	#10 counter$count = 17953;
	#10 counter$count = 17954;
	#10 counter$count = 17955;
	#10 counter$count = 17956;
	#10 counter$count = 17957;
	#10 counter$count = 17958;
	#10 counter$count = 17959;
	#10 counter$count = 17960;
	#10 counter$count = 17961;
	#10 counter$count = 17962;
	#10 counter$count = 17963;
	#10 counter$count = 17964;
	#10 counter$count = 17965;
	#10 counter$count = 17966;
	#10 counter$count = 17967;
	#10 counter$count = 17968;
	#10 counter$count = 17969;
	#10 counter$count = 17970;
	#10 counter$count = 17971;
	#10 counter$count = 17972;
	#10 counter$count = 17973;
	#10 counter$count = 17974;
	#10 counter$count = 17975;
	#10 counter$count = 17976;
	#10 counter$count = 17977;
	#10 counter$count = 17978;
	#10 counter$count = 17979;
	#10 counter$count = 17980;
	#10 counter$count = 17981;
	#10 counter$count = 17982;
	#10 counter$count = 17983;
	#10 counter$count = 17984;
	#10 counter$count = 17985;
	#10 counter$count = 17986;
	#10 counter$count = 17987;
	#10 counter$count = 17988;
	#10 counter$count = 17989;
	#10 counter$count = 17990;
	#10 counter$count = 17991;
	#10 counter$count = 17992;
	#10 counter$count = 17993;
	#10 counter$count = 17994;
	#10 counter$count = 17995;
	#10 counter$count = 17996;
	#10 counter$count = 17997;
	#10 counter$count = 17998;
	#10 counter$count = 17999;
	#10 counter$count = 18000;
	#10 counter$count = 18001;
	#10 counter$count = 18002;
	#10 counter$count = 18003;
	#10 counter$count = 18004;
	#10 counter$count = 18005;
	#10 counter$count = 18006;
	#10 counter$count = 18007;
	#10 counter$count = 18008;
	#10 counter$count = 18009;
	#10 counter$count = 18010;
	#10 counter$count = 18011;
	#10 counter$count = 18012;
	#10 counter$count = 18013;
	#10 counter$count = 18014;
	#10 counter$count = 18015;
	#10 counter$count = 18016;
	#10 counter$count = 18017;
	#10 counter$count = 18018;
	#10 counter$count = 18019;
	#10 counter$count = 18020;
	#10 counter$count = 18021;
	#10 counter$count = 18022;
	#10 counter$count = 18023;
	#10 counter$count = 18024;
	#10 counter$count = 18025;
	#10 counter$count = 18026;
	#10 counter$count = 18027;
	#10 counter$count = 18028;
	#10 counter$count = 18029;
	#10 counter$count = 18030;
	#10 counter$count = 18031;
	#10 counter$count = 18032;
	#10 counter$count = 18033;
	#10 counter$count = 18034;
	#10 counter$count = 18035;
	#10 counter$count = 18036;
	#10 counter$count = 18037;
	#10 counter$count = 18038;
	#10 counter$count = 18039;
	#10 counter$count = 18040;
	#10 counter$count = 18041;
	#10 counter$count = 18042;
	#10 counter$count = 18043;
	#10 counter$count = 18044;
	#10 counter$count = 18045;
	#10 counter$count = 18046;
	#10 counter$count = 18047;
	#10 counter$count = 18048;
	#10 counter$count = 18049;
	#10 counter$count = 18050;
	#10 counter$count = 18051;
	#10 counter$count = 18052;
	#10 counter$count = 18053;
	#10 counter$count = 18054;
	#10 counter$count = 18055;
	#10 counter$count = 18056;
	#10 counter$count = 18057;
	#10 counter$count = 18058;
	#10 counter$count = 18059;
	#10 counter$count = 18060;
	#10 counter$count = 18061;
	#10 counter$count = 18062;
	#10 counter$count = 18063;
	#10 counter$count = 18064;
	#10 counter$count = 18065;
	#10 counter$count = 18066;
	#10 counter$count = 18067;
	#10 counter$count = 18068;
	#10 counter$count = 18069;
	#10 counter$count = 18070;
	#10 counter$count = 18071;
	#10 counter$count = 18072;
	#10 counter$count = 18073;
	#10 counter$count = 18074;
	#10 counter$count = 18075;
	#10 counter$count = 18076;
	#10 counter$count = 18077;
	#10 counter$count = 18078;
	#10 counter$count = 18079;
	#10 counter$count = 18080;
	#10 counter$count = 18081;
	#10 counter$count = 18082;
	#10 counter$count = 18083;
	#10 counter$count = 18084;
	#10 counter$count = 18085;
	#10 counter$count = 18086;
	#10 counter$count = 18087;
	#10 counter$count = 18088;
	#10 counter$count = 18089;
	#10 counter$count = 18090;
	#10 counter$count = 18091;
	#10 counter$count = 18092;
	#10 counter$count = 18093;
	#10 counter$count = 18094;
	#10 counter$count = 18095;
	#10 counter$count = 18096;
	#10 counter$count = 18097;
	#10 counter$count = 18098;
	#10 counter$count = 18099;
	#10 counter$count = 18100;
	#10 counter$count = 18101;
	#10 counter$count = 18102;
	#10 counter$count = 18103;
	#10 counter$count = 18104;
	#10 counter$count = 18105;
	#10 counter$count = 18106;
	#10 counter$count = 18107;
	#10 counter$count = 18108;
	#10 counter$count = 18109;
	#10 counter$count = 18110;
	#10 counter$count = 18111;
	#10 counter$count = 18112;
	#10 counter$count = 18113;
	#10 counter$count = 18114;
	#10 counter$count = 18115;
	#10 counter$count = 18116;
	#10 counter$count = 18117;
	#10 counter$count = 18118;
	#10 counter$count = 18119;
	#10 counter$count = 18120;
	#10 counter$count = 18121;
	#10 counter$count = 18122;
	#10 counter$count = 18123;
	#10 counter$count = 18124;
	#10 counter$count = 18125;
	#10 counter$count = 18126;
	#10 counter$count = 18127;
	#10 counter$count = 18128;
	#10 counter$count = 18129;
	#10 counter$count = 18130;
	#10 counter$count = 18131;
	#10 counter$count = 18132;
	#10 counter$count = 18133;
	#10 counter$count = 18134;
	#10 counter$count = 18135;
	#10 counter$count = 18136;
	#10 counter$count = 18137;
	#10 counter$count = 18138;
	#10 counter$count = 18139;
	#10 counter$count = 18140;
	#10 counter$count = 18141;
	#10 counter$count = 18142;
	#10 counter$count = 18143;
	#10 counter$count = 18144;
	#10 counter$count = 18145;
	#10 counter$count = 18146;
	#10 counter$count = 18147;
	#10 counter$count = 18148;
	#10 counter$count = 18149;
	#10 counter$count = 18150;
	#10 counter$count = 18151;
	#10 counter$count = 18152;
	#10 counter$count = 18153;
	#10 counter$count = 18154;
	#10 counter$count = 18155;
	#10 counter$count = 18156;
	#10 counter$count = 18157;
	#10 counter$count = 18158;
	#10 counter$count = 18159;
	#10 counter$count = 18160;
	#10 counter$count = 18161;
	#10 counter$count = 18162;
	#10 counter$count = 18163;
	#10 counter$count = 18164;
	#10 counter$count = 18165;
	#10 counter$count = 18166;
	#10 counter$count = 18167;
	#10 counter$count = 18168;
	#10 counter$count = 18169;
	#10 counter$count = 18170;
	#10 counter$count = 18171;
	#10 counter$count = 18172;
	#10 counter$count = 18173;
	#10 counter$count = 18174;
	#10 counter$count = 18175;
	#10 counter$count = 18176;
	#10 counter$count = 18177;
	#10 counter$count = 18178;
	#10 counter$count = 18179;
	#10 counter$count = 18180;
	#10 counter$count = 18181;
	#10 counter$count = 18182;
	#10 counter$count = 18183;
	#10 counter$count = 18184;
	#10 counter$count = 18185;
	#10 counter$count = 18186;
	#10 counter$count = 18187;
	#10 counter$count = 18188;
	#10 counter$count = 18189;
	#10 counter$count = 18190;
	#10 counter$count = 18191;
	#10 counter$count = 18192;
	#10 counter$count = 18193;
	#10 counter$count = 18194;
	#10 counter$count = 18195;
	#10 counter$count = 18196;
	#10 counter$count = 18197;
	#10 counter$count = 18198;
	#10 counter$count = 18199;
	#10 counter$count = 18200;
	#10 counter$count = 18201;
	#10 counter$count = 18202;
	#10 counter$count = 18203;
	#10 counter$count = 18204;
	#10 counter$count = 18205;
	#10 counter$count = 18206;
	#10 counter$count = 18207;
	#10 counter$count = 18208;
	#10 counter$count = 18209;
	#10 counter$count = 18210;
	#10 counter$count = 18211;
	#10 counter$count = 18212;
	#10 counter$count = 18213;
	#10 counter$count = 18214;
	#10 counter$count = 18215;
	#10 counter$count = 18216;
	#10 counter$count = 18217;
	#10 counter$count = 18218;
	#10 counter$count = 18219;
	#10 counter$count = 18220;
	#10 counter$count = 18221;
	#10 counter$count = 18222;
	#10 counter$count = 18223;
	#10 counter$count = 18224;
	#10 counter$count = 18225;
	#10 counter$count = 18226;
	#10 counter$count = 18227;
	#10 counter$count = 18228;
	#10 counter$count = 18229;
	#10 counter$count = 18230;
	#10 counter$count = 18231;
	#10 counter$count = 18232;
	#10 counter$count = 18233;
	#10 counter$count = 18234;
	#10 counter$count = 18235;
	#10 counter$count = 18236;
	#10 counter$count = 18237;
	#10 counter$count = 18238;
	#10 counter$count = 18239;
	#10 counter$count = 18240;
	#10 counter$count = 18241;
	#10 counter$count = 18242;
	#10 counter$count = 18243;
	#10 counter$count = 18244;
	#10 counter$count = 18245;
	#10 counter$count = 18246;
	#10 counter$count = 18247;
	#10 counter$count = 18248;
	#10 counter$count = 18249;
	#10 counter$count = 18250;
	#10 counter$count = 18251;
	#10 counter$count = 18252;
	#10 counter$count = 18253;
	#10 counter$count = 18254;
	#10 counter$count = 18255;
	#10 counter$count = 18256;
	#10 counter$count = 18257;
	#10 counter$count = 18258;
	#10 counter$count = 18259;
	#10 counter$count = 18260;
	#10 counter$count = 18261;
	#10 counter$count = 18262;
	#10 counter$count = 18263;
	#10 counter$count = 18264;
	#10 counter$count = 18265;
	#10 counter$count = 18266;
	#10 counter$count = 18267;
	#10 counter$count = 18268;
	#10 counter$count = 18269;
	#10 counter$count = 18270;
	#10 counter$count = 18271;
	#10 counter$count = 18272;
	#10 counter$count = 18273;
	#10 counter$count = 18274;
	#10 counter$count = 18275;
	#10 counter$count = 18276;
	#10 counter$count = 18277;
	#10 counter$count = 18278;
	#10 counter$count = 18279;
	#10 counter$count = 18280;
	#10 counter$count = 18281;
	#10 counter$count = 18282;
	#10 counter$count = 18283;
	#10 counter$count = 18284;
	#10 counter$count = 18285;
	#10 counter$count = 18286;
	#10 counter$count = 18287;
	#10 counter$count = 18288;
	#10 counter$count = 18289;
	#10 counter$count = 18290;
	#10 counter$count = 18291;
	#10 counter$count = 18292;
	#10 counter$count = 18293;
	#10 counter$count = 18294;
	#10 counter$count = 18295;
	#10 counter$count = 18296;
	#10 counter$count = 18297;
	#10 counter$count = 18298;
	#10 counter$count = 18299;
	#10 counter$count = 18300;
	#10 counter$count = 18301;
	#10 counter$count = 18302;
	#10 counter$count = 18303;
	#10 counter$count = 18304;
	#10 counter$count = 18305;
	#10 counter$count = 18306;
	#10 counter$count = 18307;
	#10 counter$count = 18308;
	#10 counter$count = 18309;
	#10 counter$count = 18310;
	#10 counter$count = 18311;
	#10 counter$count = 18312;
	#10 counter$count = 18313;
	#10 counter$count = 18314;
	#10 counter$count = 18315;
	#10 counter$count = 18316;
	#10 counter$count = 18317;
	#10 counter$count = 18318;
	#10 counter$count = 18319;
	#10 counter$count = 18320;
	#10 counter$count = 18321;
	#10 counter$count = 18322;
	#10 counter$count = 18323;
	#10 counter$count = 18324;
	#10 counter$count = 18325;
	#10 counter$count = 18326;
	#10 counter$count = 18327;
	#10 counter$count = 18328;
	#10 counter$count = 18329;
	#10 counter$count = 18330;
	#10 counter$count = 18331;
	#10 counter$count = 18332;
	#10 counter$count = 18333;
	#10 counter$count = 18334;
	#10 counter$count = 18335;
	#10 counter$count = 18336;
	#10 counter$count = 18337;
	#10 counter$count = 18338;
	#10 counter$count = 18339;
	#10 counter$count = 18340;
	#10 counter$count = 18341;
	#10 counter$count = 18342;
	#10 counter$count = 18343;
	#10 counter$count = 18344;
	#10 counter$count = 18345;
	#10 counter$count = 18346;
	#10 counter$count = 18347;
	#10 counter$count = 18348;
	#10 counter$count = 18349;
	#10 counter$count = 18350;
	#10 counter$count = 18351;
	#10 counter$count = 18352;
	#10 counter$count = 18353;
	#10 counter$count = 18354;
	#10 counter$count = 18355;
	#10 counter$count = 18356;
	#10 counter$count = 18357;
	#10 counter$count = 18358;
	#10 counter$count = 18359;
	#10 counter$count = 18360;
	#10 counter$count = 18361;
	#10 counter$count = 18362;
	#10 counter$count = 18363;
	#10 counter$count = 18364;
	#10 counter$count = 18365;
	#10 counter$count = 18366;
	#10 counter$count = 18367;
	#10 counter$count = 18368;
	#10 counter$count = 18369;
	#10 counter$count = 18370;
	#10 counter$count = 18371;
	#10 counter$count = 18372;
	#10 counter$count = 18373;
	#10 counter$count = 18374;
	#10 counter$count = 18375;
	#10 counter$count = 18376;
	#10 counter$count = 18377;
	#10 counter$count = 18378;
	#10 counter$count = 18379;
	#10 counter$count = 18380;
	#10 counter$count = 18381;
	#10 counter$count = 18382;
	#10 counter$count = 18383;
	#10 counter$count = 18384;
	#10 counter$count = 18385;
	#10 counter$count = 18386;
	#10 counter$count = 18387;
	#10 counter$count = 18388;
	#10 counter$count = 18389;
	#10 counter$count = 18390;
	#10 counter$count = 18391;
	#10 counter$count = 18392;
	#10 counter$count = 18393;
	#10 counter$count = 18394;
	#10 counter$count = 18395;
	#10 counter$count = 18396;
	#10 counter$count = 18397;
	#10 counter$count = 18398;
	#10 counter$count = 18399;
	#10 counter$count = 18400;
	#10 counter$count = 18401;
	#10 counter$count = 18402;
	#10 counter$count = 18403;
	#10 counter$count = 18404;
	#10 counter$count = 18405;
	#10 counter$count = 18406;
	#10 counter$count = 18407;
	#10 counter$count = 18408;
	#10 counter$count = 18409;
	#10 counter$count = 18410;
	#10 counter$count = 18411;
	#10 counter$count = 18412;
	#10 counter$count = 18413;
	#10 counter$count = 18414;
	#10 counter$count = 18415;
	#10 counter$count = 18416;
	#10 counter$count = 18417;
	#10 counter$count = 18418;
	#10 counter$count = 18419;
	#10 counter$count = 18420;
	#10 counter$count = 18421;
	#10 counter$count = 18422;
	#10 counter$count = 18423;
	#10 counter$count = 18424;
	#10 counter$count = 18425;
	#10 counter$count = 18426;
	#10 counter$count = 18427;
	#10 counter$count = 18428;
	#10 counter$count = 18429;
	#10 counter$count = 18430;
	#10 counter$count = 18431;
	#10 counter$count = 18432;
	#10 counter$count = 18433;
	#10 counter$count = 18434;
	#10 counter$count = 18435;
	#10 counter$count = 18436;
	#10 counter$count = 18437;
	#10 counter$count = 18438;
	#10 counter$count = 18439;
	#10 counter$count = 18440;
	#10 counter$count = 18441;
	#10 counter$count = 18442;
	#10 counter$count = 18443;
	#10 counter$count = 18444;
	#10 counter$count = 18445;
	#10 counter$count = 18446;
	#10 counter$count = 18447;
	#10 counter$count = 18448;
	#10 counter$count = 18449;
	#10 counter$count = 18450;
	#10 counter$count = 18451;
	#10 counter$count = 18452;
	#10 counter$count = 18453;
	#10 counter$count = 18454;
	#10 counter$count = 18455;
	#10 counter$count = 18456;
	#10 counter$count = 18457;
	#10 counter$count = 18458;
	#10 counter$count = 18459;
	#10 counter$count = 18460;
	#10 counter$count = 18461;
	#10 counter$count = 18462;
	#10 counter$count = 18463;
	#10 counter$count = 18464;
	#10 counter$count = 18465;
	#10 counter$count = 18466;
	#10 counter$count = 18467;
	#10 counter$count = 18468;
	#10 counter$count = 18469;
	#10 counter$count = 18470;
	#10 counter$count = 18471;
	#10 counter$count = 18472;
	#10 counter$count = 18473;
	#10 counter$count = 18474;
	#10 counter$count = 18475;
	#10 counter$count = 18476;
	#10 counter$count = 18477;
	#10 counter$count = 18478;
	#10 counter$count = 18479;
	#10 counter$count = 18480;
	#10 counter$count = 18481;
	#10 counter$count = 18482;
	#10 counter$count = 18483;
	#10 counter$count = 18484;
	#10 counter$count = 18485;
	#10 counter$count = 18486;
	#10 counter$count = 18487;
	#10 counter$count = 18488;
	#10 counter$count = 18489;
	#10 counter$count = 18490;
	#10 counter$count = 18491;
	#10 counter$count = 18492;
	#10 counter$count = 18493;
	#10 counter$count = 18494;
	#10 counter$count = 18495;
	#10 counter$count = 18496;
	#10 counter$count = 18497;
	#10 counter$count = 18498;
	#10 counter$count = 18499;
	#10 counter$count = 18500;
	#10 counter$count = 18501;
	#10 counter$count = 18502;
	#10 counter$count = 18503;
	#10 counter$count = 18504;
	#10 counter$count = 18505;
	#10 counter$count = 18506;
	#10 counter$count = 18507;
	#10 counter$count = 18508;
	#10 counter$count = 18509;
	#10 counter$count = 18510;
	#10 counter$count = 18511;
	#10 counter$count = 18512;
	#10 counter$count = 18513;
	#10 counter$count = 18514;
	#10 counter$count = 18515;
	#10 counter$count = 18516;
	#10 counter$count = 18517;
	#10 counter$count = 18518;
	#10 counter$count = 18519;
	#10 counter$count = 18520;
	#10 counter$count = 18521;
	#10 counter$count = 18522;
	#10 counter$count = 18523;
	#10 counter$count = 18524;
	#10 counter$count = 18525;
	#10 counter$count = 18526;
	#10 counter$count = 18527;
	#10 counter$count = 18528;
	#10 counter$count = 18529;
	#10 counter$count = 18530;
	#10 counter$count = 18531;
	#10 counter$count = 18532;
	#10 counter$count = 18533;
	#10 counter$count = 18534;
	#10 counter$count = 18535;
	#10 counter$count = 18536;
	#10 counter$count = 18537;
	#10 counter$count = 18538;
	#10 counter$count = 18539;
	#10 counter$count = 18540;
	#10 counter$count = 18541;
	#10 counter$count = 18542;
	#10 counter$count = 18543;
	#10 counter$count = 18544;
	#10 counter$count = 18545;
	#10 counter$count = 18546;
	#10 counter$count = 18547;
	#10 counter$count = 18548;
	#10 counter$count = 18549;
	#10 counter$count = 18550;
	#10 counter$count = 18551;
	#10 counter$count = 18552;
	#10 counter$count = 18553;
	#10 counter$count = 18554;
	#10 counter$count = 18555;
	#10 counter$count = 18556;
	#10 counter$count = 18557;
	#10 counter$count = 18558;
	#10 counter$count = 18559;
	#10 counter$count = 18560;
	#10 counter$count = 18561;
	#10 counter$count = 18562;
	#10 counter$count = 18563;
	#10 counter$count = 18564;
	#10 counter$count = 18565;
	#10 counter$count = 18566;
	#10 counter$count = 18567;
	#10 counter$count = 18568;
	#10 counter$count = 18569;
	#10 counter$count = 18570;
	#10 counter$count = 18571;
	#10 counter$count = 18572;
	#10 counter$count = 18573;
	#10 counter$count = 18574;
	#10 counter$count = 18575;
	#10 counter$count = 18576;
	#10 counter$count = 18577;
	#10 counter$count = 18578;
	#10 counter$count = 18579;
	#10 counter$count = 18580;
	#10 counter$count = 18581;
	#10 counter$count = 18582;
	#10 counter$count = 18583;
	#10 counter$count = 18584;
	#10 counter$count = 18585;
	#10 counter$count = 18586;
	#10 counter$count = 18587;
	#10 counter$count = 18588;
	#10 counter$count = 18589;
	#10 counter$count = 18590;
	#10 counter$count = 18591;
	#10 counter$count = 18592;
	#10 counter$count = 18593;
	#10 counter$count = 18594;
	#10 counter$count = 18595;
	#10 counter$count = 18596;
	#10 counter$count = 18597;
	#10 counter$count = 18598;
	#10 counter$count = 18599;
	#10 counter$count = 18600;
	#10 counter$count = 18601;
	#10 counter$count = 18602;
	#10 counter$count = 18603;
	#10 counter$count = 18604;
	#10 counter$count = 18605;
	#10 counter$count = 18606;
	#10 counter$count = 18607;
	#10 counter$count = 18608;
	#10 counter$count = 18609;
	#10 counter$count = 18610;
	#10 counter$count = 18611;
	#10 counter$count = 18612;
	#10 counter$count = 18613;
	#10 counter$count = 18614;
	#10 counter$count = 18615;
	#10 counter$count = 18616;
	#10 counter$count = 18617;
	#10 counter$count = 18618;
	#10 counter$count = 18619;
	#10 counter$count = 18620;
	#10 counter$count = 18621;
	#10 counter$count = 18622;
	#10 counter$count = 18623;
	#10 counter$count = 18624;
	#10 counter$count = 18625;
	#10 counter$count = 18626;
	#10 counter$count = 18627;
	#10 counter$count = 18628;
	#10 counter$count = 18629;
	#10 counter$count = 18630;
	#10 counter$count = 18631;
	#10 counter$count = 18632;
	#10 counter$count = 18633;
	#10 counter$count = 18634;
	#10 counter$count = 18635;
	#10 counter$count = 18636;
	#10 counter$count = 18637;
	#10 counter$count = 18638;
	#10 counter$count = 18639;
	#10 counter$count = 18640;
	#10 counter$count = 18641;
	#10 counter$count = 18642;
	#10 counter$count = 18643;
	#10 counter$count = 18644;
	#10 counter$count = 18645;
	#10 counter$count = 18646;
	#10 counter$count = 18647;
	#10 counter$count = 18648;
	#10 counter$count = 18649;
	#10 counter$count = 18650;
	#10 counter$count = 18651;
	#10 counter$count = 18652;
	#10 counter$count = 18653;
	#10 counter$count = 18654;
	#10 counter$count = 18655;
	#10 counter$count = 18656;
	#10 counter$count = 18657;
	#10 counter$count = 18658;
	#10 counter$count = 18659;
	#10 counter$count = 18660;
	#10 counter$count = 18661;
	#10 counter$count = 18662;
	#10 counter$count = 18663;
	#10 counter$count = 18664;
	#10 counter$count = 18665;
	#10 counter$count = 18666;
	#10 counter$count = 18667;
	#10 counter$count = 18668;
	#10 counter$count = 18669;
	#10 counter$count = 18670;
	#10 counter$count = 18671;
	#10 counter$count = 18672;
	#10 counter$count = 18673;
	#10 counter$count = 18674;
	#10 counter$count = 18675;
	#10 counter$count = 18676;
	#10 counter$count = 18677;
	#10 counter$count = 18678;
	#10 counter$count = 18679;
	#10 counter$count = 18680;
	#10 counter$count = 18681;
	#10 counter$count = 18682;
	#10 counter$count = 18683;
	#10 counter$count = 18684;
	#10 counter$count = 18685;
	#10 counter$count = 18686;
	#10 counter$count = 18687;
	#10 counter$count = 18688;
	#10 counter$count = 18689;
	#10 counter$count = 18690;
	#10 counter$count = 18691;
	#10 counter$count = 18692;
	#10 counter$count = 18693;
	#10 counter$count = 18694;
	#10 counter$count = 18695;
	#10 counter$count = 18696;
	#10 counter$count = 18697;
	#10 counter$count = 18698;
	#10 counter$count = 18699;
	#10 counter$count = 18700;
	#10 counter$count = 18701;
	#10 counter$count = 18702;
	#10 counter$count = 18703;
	#10 counter$count = 18704;
	#10 counter$count = 18705;
	#10 counter$count = 18706;
	#10 counter$count = 18707;
	#10 counter$count = 18708;
	#10 counter$count = 18709;
	#10 counter$count = 18710;
	#10 counter$count = 18711;
	#10 counter$count = 18712;
	#10 counter$count = 18713;
	#10 counter$count = 18714;
	#10 counter$count = 18715;
	#10 counter$count = 18716;
	#10 counter$count = 18717;
	#10 counter$count = 18718;
	#10 counter$count = 18719;
	#10 counter$count = 18720;
	#10 counter$count = 18721;
	#10 counter$count = 18722;
	#10 counter$count = 18723;
	#10 counter$count = 18724;
	#10 counter$count = 18725;
	#10 counter$count = 18726;
	#10 counter$count = 18727;
	#10 counter$count = 18728;
	#10 counter$count = 18729;
	#10 counter$count = 18730;
	#10 counter$count = 18731;
	#10 counter$count = 18732;
	#10 counter$count = 18733;
	#10 counter$count = 18734;
	#10 counter$count = 18735;
	#10 counter$count = 18736;
	#10 counter$count = 18737;
	#10 counter$count = 18738;
	#10 counter$count = 18739;
	#10 counter$count = 18740;
	#10 counter$count = 18741;
	#10 counter$count = 18742;
	#10 counter$count = 18743;
	#10 counter$count = 18744;
	#10 counter$count = 18745;
	#10 counter$count = 18746;
	#10 counter$count = 18747;
	#10 counter$count = 18748;
	#10 counter$count = 18749;
	#10 counter$count = 18750;
	#10 counter$count = 18751;
	#10 counter$count = 18752;
	#10 counter$count = 18753;
	#10 counter$count = 18754;
	#10 counter$count = 18755;
	#10 counter$count = 18756;
	#10 counter$count = 18757;
	#10 counter$count = 18758;
	#10 counter$count = 18759;
	#10 counter$count = 18760;
	#10 counter$count = 18761;
	#10 counter$count = 18762;
	#10 counter$count = 18763;
	#10 counter$count = 18764;
	#10 counter$count = 18765;
	#10 counter$count = 18766;
	#10 counter$count = 18767;
	#10 counter$count = 18768;
	#10 counter$count = 18769;
	#10 counter$count = 18770;
	#10 counter$count = 18771;
	#10 counter$count = 18772;
	#10 counter$count = 18773;
	#10 counter$count = 18774;
	#10 counter$count = 18775;
	#10 counter$count = 18776;
	#10 counter$count = 18777;
	#10 counter$count = 18778;
	#10 counter$count = 18779;
	#10 counter$count = 18780;
	#10 counter$count = 18781;
	#10 counter$count = 18782;
	#10 counter$count = 18783;
	#10 counter$count = 18784;
	#10 counter$count = 18785;
	#10 counter$count = 18786;
	#10 counter$count = 18787;
	#10 counter$count = 18788;
	#10 counter$count = 18789;
	#10 counter$count = 18790;
	#10 counter$count = 18791;
	#10 counter$count = 18792;
	#10 counter$count = 18793;
	#10 counter$count = 18794;
	#10 counter$count = 18795;
	#10 counter$count = 18796;
	#10 counter$count = 18797;
	#10 counter$count = 18798;
	#10 counter$count = 18799;
	#10 counter$count = 18800;
	#10 counter$count = 18801;
	#10 counter$count = 18802;
	#10 counter$count = 18803;
	#10 counter$count = 18804;
	#10 counter$count = 18805;
	#10 counter$count = 18806;
	#10 counter$count = 18807;
	#10 counter$count = 18808;
	#10 counter$count = 18809;
	#10 counter$count = 18810;
	#10 counter$count = 18811;
	#10 counter$count = 18812;
	#10 counter$count = 18813;
	#10 counter$count = 18814;
	#10 counter$count = 18815;
	#10 counter$count = 18816;
	#10 counter$count = 18817;
	#10 counter$count = 18818;
	#10 counter$count = 18819;
	#10 counter$count = 18820;
	#10 counter$count = 18821;
	#10 counter$count = 18822;
	#10 counter$count = 18823;
	#10 counter$count = 18824;
	#10 counter$count = 18825;
	#10 counter$count = 18826;
	#10 counter$count = 18827;
	#10 counter$count = 18828;
	#10 counter$count = 18829;
	#10 counter$count = 18830;
	#10 counter$count = 18831;
	#10 counter$count = 18832;
	#10 counter$count = 18833;
	#10 counter$count = 18834;
	#10 counter$count = 18835;
	#10 counter$count = 18836;
	#10 counter$count = 18837;
	#10 counter$count = 18838;
	#10 counter$count = 18839;
	#10 counter$count = 18840;
	#10 counter$count = 18841;
	#10 counter$count = 18842;
	#10 counter$count = 18843;
	#10 counter$count = 18844;
	#10 counter$count = 18845;
	#10 counter$count = 18846;
	#10 counter$count = 18847;
	#10 counter$count = 18848;
	#10 counter$count = 18849;
	#10 counter$count = 18850;
	#10 counter$count = 18851;
	#10 counter$count = 18852;
	#10 counter$count = 18853;
	#10 counter$count = 18854;
	#10 counter$count = 18855;
	#10 counter$count = 18856;
	#10 counter$count = 18857;
	#10 counter$count = 18858;
	#10 counter$count = 18859;
	#10 counter$count = 18860;
	#10 counter$count = 18861;
	#10 counter$count = 18862;
	#10 counter$count = 18863;
	#10 counter$count = 18864;
	#10 counter$count = 18865;
	#10 counter$count = 18866;
	#10 counter$count = 18867;
	#10 counter$count = 18868;
	#10 counter$count = 18869;
	#10 counter$count = 18870;
	#10 counter$count = 18871;
	#10 counter$count = 18872;
	#10 counter$count = 18873;
	#10 counter$count = 18874;
	#10 counter$count = 18875;
	#10 counter$count = 18876;
	#10 counter$count = 18877;
	#10 counter$count = 18878;
	#10 counter$count = 18879;
	#10 counter$count = 18880;
	#10 counter$count = 18881;
	#10 counter$count = 18882;
	#10 counter$count = 18883;
	#10 counter$count = 18884;
	#10 counter$count = 18885;
	#10 counter$count = 18886;
	#10 counter$count = 18887;
	#10 counter$count = 18888;
	#10 counter$count = 18889;
	#10 counter$count = 18890;
	#10 counter$count = 18891;
	#10 counter$count = 18892;
	#10 counter$count = 18893;
	#10 counter$count = 18894;
	#10 counter$count = 18895;
	#10 counter$count = 18896;
	#10 counter$count = 18897;
	#10 counter$count = 18898;
	#10 counter$count = 18899;
	#10 counter$count = 18900;
	#10 counter$count = 18901;
	#10 counter$count = 18902;
	#10 counter$count = 18903;
	#10 counter$count = 18904;
	#10 counter$count = 18905;
	#10 counter$count = 18906;
	#10 counter$count = 18907;
	#10 counter$count = 18908;
	#10 counter$count = 18909;
	#10 counter$count = 18910;
	#10 counter$count = 18911;
	#10 counter$count = 18912;
	#10 counter$count = 18913;
	#10 counter$count = 18914;
	#10 counter$count = 18915;
	#10 counter$count = 18916;
	#10 counter$count = 18917;
	#10 counter$count = 18918;
	#10 counter$count = 18919;
	#10 counter$count = 18920;
	#10 counter$count = 18921;
	#10 counter$count = 18922;
	#10 counter$count = 18923;
	#10 counter$count = 18924;
	#10 counter$count = 18925;
	#10 counter$count = 18926;
	#10 counter$count = 18927;
	#10 counter$count = 18928;
	#10 counter$count = 18929;
	#10 counter$count = 18930;
	#10 counter$count = 18931;
	#10 counter$count = 18932;
	#10 counter$count = 18933;
	#10 counter$count = 18934;
	#10 counter$count = 18935;
	#10 counter$count = 18936;
	#10 counter$count = 18937;
	#10 counter$count = 18938;
	#10 counter$count = 18939;
	#10 counter$count = 18940;
	#10 counter$count = 18941;
	#10 counter$count = 18942;
	#10 counter$count = 18943;
	#10 counter$count = 18944;
	#10 counter$count = 18945;
	#10 counter$count = 18946;
	#10 counter$count = 18947;
	#10 counter$count = 18948;
	#10 counter$count = 18949;
	#10 counter$count = 18950;
	#10 counter$count = 18951;
	#10 counter$count = 18952;
	#10 counter$count = 18953;
	#10 counter$count = 18954;
	#10 counter$count = 18955;
	#10 counter$count = 18956;
	#10 counter$count = 18957;
	#10 counter$count = 18958;
	#10 counter$count = 18959;
	#10 counter$count = 18960;
	#10 counter$count = 18961;
	#10 counter$count = 18962;
	#10 counter$count = 18963;
	#10 counter$count = 18964;
	#10 counter$count = 18965;
	#10 counter$count = 18966;
	#10 counter$count = 18967;
	#10 counter$count = 18968;
	#10 counter$count = 18969;
	#10 counter$count = 18970;
	#10 counter$count = 18971;
	#10 counter$count = 18972;
	#10 counter$count = 18973;
	#10 counter$count = 18974;
	#10 counter$count = 18975;
	#10 counter$count = 18976;
	#10 counter$count = 18977;
	#10 counter$count = 18978;
	#10 counter$count = 18979;
	#10 counter$count = 18980;
	#10 counter$count = 18981;
	#10 counter$count = 18982;
	#10 counter$count = 18983;
	#10 counter$count = 18984;
	#10 counter$count = 18985;
	#10 counter$count = 18986;
	#10 counter$count = 18987;
	#10 counter$count = 18988;
	#10 counter$count = 18989;
	#10 counter$count = 18990;
	#10 counter$count = 18991;
	#10 counter$count = 18992;
	#10 counter$count = 18993;
	#10 counter$count = 18994;
	#10 counter$count = 18995;
	#10 counter$count = 18996;
	#10 counter$count = 18997;
	#10 counter$count = 18998;
	#10 counter$count = 18999;
	#10 counter$count = 19000;
	#10 counter$count = 19001;
	#10 counter$count = 19002;
	#10 counter$count = 19003;
	#10 counter$count = 19004;
	#10 counter$count = 19005;
	#10 counter$count = 19006;
	#10 counter$count = 19007;
	#10 counter$count = 19008;
	#10 counter$count = 19009;
	#10 counter$count = 19010;
	#10 counter$count = 19011;
	#10 counter$count = 19012;
	#10 counter$count = 19013;
	#10 counter$count = 19014;
	#10 counter$count = 19015;
	#10 counter$count = 19016;
	#10 counter$count = 19017;
	#10 counter$count = 19018;
	#10 counter$count = 19019;
	#10 counter$count = 19020;
	#10 counter$count = 19021;
	#10 counter$count = 19022;
	#10 counter$count = 19023;
	#10 counter$count = 19024;
	#10 counter$count = 19025;
	#10 counter$count = 19026;
	#10 counter$count = 19027;
	#10 counter$count = 19028;
	#10 counter$count = 19029;
	#10 counter$count = 19030;
	#10 counter$count = 19031;
	#10 counter$count = 19032;
	#10 counter$count = 19033;
	#10 counter$count = 19034;
	#10 counter$count = 19035;
	#10 counter$count = 19036;
	#10 counter$count = 19037;
	#10 counter$count = 19038;
	#10 counter$count = 19039;
	#10 counter$count = 19040;
	#10 counter$count = 19041;
	#10 counter$count = 19042;
	#10 counter$count = 19043;
	#10 counter$count = 19044;
	#10 counter$count = 19045;
	#10 counter$count = 19046;
	#10 counter$count = 19047;
	#10 counter$count = 19048;
	#10 counter$count = 19049;
	#10 counter$count = 19050;
	#10 counter$count = 19051;
	#10 counter$count = 19052;
	#10 counter$count = 19053;
	#10 counter$count = 19054;
	#10 counter$count = 19055;
	#10 counter$count = 19056;
	#10 counter$count = 19057;
	#10 counter$count = 19058;
	#10 counter$count = 19059;
	#10 counter$count = 19060;
	#10 counter$count = 19061;
	#10 counter$count = 19062;
	#10 counter$count = 19063;
	#10 counter$count = 19064;
	#10 counter$count = 19065;
	#10 counter$count = 19066;
	#10 counter$count = 19067;
	#10 counter$count = 19068;
	#10 counter$count = 19069;
	#10 counter$count = 19070;
	#10 counter$count = 19071;
	#10 counter$count = 19072;
	#10 counter$count = 19073;
	#10 counter$count = 19074;
	#10 counter$count = 19075;
	#10 counter$count = 19076;
	#10 counter$count = 19077;
	#10 counter$count = 19078;
	#10 counter$count = 19079;
	#10 counter$count = 19080;
	#10 counter$count = 19081;
	#10 counter$count = 19082;
	#10 counter$count = 19083;
	#10 counter$count = 19084;
	#10 counter$count = 19085;
	#10 counter$count = 19086;
	#10 counter$count = 19087;
	#10 counter$count = 19088;
	#10 counter$count = 19089;
	#10 counter$count = 19090;
	#10 counter$count = 19091;
	#10 counter$count = 19092;
	#10 counter$count = 19093;
	#10 counter$count = 19094;
	#10 counter$count = 19095;
	#10 counter$count = 19096;
	#10 counter$count = 19097;
	#10 counter$count = 19098;
	#10 counter$count = 19099;
	#10 counter$count = 19100;
	#10 counter$count = 19101;
	#10 counter$count = 19102;
	#10 counter$count = 19103;
	#10 counter$count = 19104;
	#10 counter$count = 19105;
	#10 counter$count = 19106;
	#10 counter$count = 19107;
	#10 counter$count = 19108;
	#10 counter$count = 19109;
	#10 counter$count = 19110;
	#10 counter$count = 19111;
	#10 counter$count = 19112;
	#10 counter$count = 19113;
	#10 counter$count = 19114;
	#10 counter$count = 19115;
	#10 counter$count = 19116;
	#10 counter$count = 19117;
	#10 counter$count = 19118;
	#10 counter$count = 19119;
	#10 counter$count = 19120;
	#10 counter$count = 19121;
	#10 counter$count = 19122;
	#10 counter$count = 19123;
	#10 counter$count = 19124;
	#10 counter$count = 19125;
	#10 counter$count = 19126;
	#10 counter$count = 19127;
	#10 counter$count = 19128;
	#10 counter$count = 19129;
	#10 counter$count = 19130;
	#10 counter$count = 19131;
	#10 counter$count = 19132;
	#10 counter$count = 19133;
	#10 counter$count = 19134;
	#10 counter$count = 19135;
	#10 counter$count = 19136;
	#10 counter$count = 19137;
	#10 counter$count = 19138;
	#10 counter$count = 19139;
	#10 counter$count = 19140;
	#10 counter$count = 19141;
	#10 counter$count = 19142;
	#10 counter$count = 19143;
	#10 counter$count = 19144;
	#10 counter$count = 19145;
	#10 counter$count = 19146;
	#10 counter$count = 19147;
	#10 counter$count = 19148;
	#10 counter$count = 19149;
	#10 counter$count = 19150;
	#10 counter$count = 19151;
	#10 counter$count = 19152;
	#10 counter$count = 19153;
	#10 counter$count = 19154;
	#10 counter$count = 19155;
	#10 counter$count = 19156;
	#10 counter$count = 19157;
	#10 counter$count = 19158;
	#10 counter$count = 19159;
	#10 counter$count = 19160;
	#10 counter$count = 19161;
	#10 counter$count = 19162;
	#10 counter$count = 19163;
	#10 counter$count = 19164;
	#10 counter$count = 19165;
	#10 counter$count = 19166;
	#10 counter$count = 19167;
	#10 counter$count = 19168;
	#10 counter$count = 19169;
	#10 counter$count = 19170;
	#10 counter$count = 19171;
	#10 counter$count = 19172;
	#10 counter$count = 19173;
	#10 counter$count = 19174;
	#10 counter$count = 19175;
	#10 counter$count = 19176;
	#10 counter$count = 19177;
	#10 counter$count = 19178;
	#10 counter$count = 19179;
	#10 counter$count = 19180;
	#10 counter$count = 19181;
	#10 counter$count = 19182;
	#10 counter$count = 19183;
	#10 counter$count = 19184;
	#10 counter$count = 19185;
	#10 counter$count = 19186;
	#10 counter$count = 19187;
	#10 counter$count = 19188;
	#10 counter$count = 19189;
	#10 counter$count = 19190;
	#10 counter$count = 19191;
	#10 counter$count = 19192;
	#10 counter$count = 19193;
	#10 counter$count = 19194;
	#10 counter$count = 19195;
	#10 counter$count = 19196;
	#10 counter$count = 19197;
	#10 counter$count = 19198;
	#10 counter$count = 19199;
	#10 counter$count = 19200;
	#10 counter$count = 19201;
	#10 counter$count = 19202;
	#10 counter$count = 19203;
	#10 counter$count = 19204;
	#10 counter$count = 19205;
	#10 counter$count = 19206;
	#10 counter$count = 19207;
	#10 counter$count = 19208;
	#10 counter$count = 19209;
	#10 counter$count = 19210;
	#10 counter$count = 19211;
	#10 counter$count = 19212;
	#10 counter$count = 19213;
	#10 counter$count = 19214;
	#10 counter$count = 19215;
	#10 counter$count = 19216;
	#10 counter$count = 19217;
	#10 counter$count = 19218;
	#10 counter$count = 19219;
	#10 counter$count = 19220;
	#10 counter$count = 19221;
	#10 counter$count = 19222;
	#10 counter$count = 19223;
	#10 counter$count = 19224;
	#10 counter$count = 19225;
	#10 counter$count = 19226;
	#10 counter$count = 19227;
	#10 counter$count = 19228;
	#10 counter$count = 19229;
	#10 counter$count = 19230;
	#10 counter$count = 19231;
	#10 counter$count = 19232;
	#10 counter$count = 19233;
	#10 counter$count = 19234;
	#10 counter$count = 19235;
	#10 counter$count = 19236;
	#10 counter$count = 19237;
	#10 counter$count = 19238;
	#10 counter$count = 19239;
	#10 counter$count = 19240;
	#10 counter$count = 19241;
	#10 counter$count = 19242;
	#10 counter$count = 19243;
	#10 counter$count = 19244;
	#10 counter$count = 19245;
	#10 counter$count = 19246;
	#10 counter$count = 19247;
	#10 counter$count = 19248;
	#10 counter$count = 19249;
	#10 counter$count = 19250;
	#10 counter$count = 19251;
	#10 counter$count = 19252;
	#10 counter$count = 19253;
	#10 counter$count = 19254;
	#10 counter$count = 19255;
	#10 counter$count = 19256;
	#10 counter$count = 19257;
	#10 counter$count = 19258;
	#10 counter$count = 19259;
	#10 counter$count = 19260;
	#10 counter$count = 19261;
	#10 counter$count = 19262;
	#10 counter$count = 19263;
	#10 counter$count = 19264;
	#10 counter$count = 19265;
	#10 counter$count = 19266;
	#10 counter$count = 19267;
	#10 counter$count = 19268;
	#10 counter$count = 19269;
	#10 counter$count = 19270;
	#10 counter$count = 19271;
	#10 counter$count = 19272;
	#10 counter$count = 19273;
	#10 counter$count = 19274;
	#10 counter$count = 19275;
	#10 counter$count = 19276;
	#10 counter$count = 19277;
	#10 counter$count = 19278;
	#10 counter$count = 19279;
	#10 counter$count = 19280;
	#10 counter$count = 19281;
	#10 counter$count = 19282;
	#10 counter$count = 19283;
	#10 counter$count = 19284;
	#10 counter$count = 19285;
	#10 counter$count = 19286;
	#10 counter$count = 19287;
	#10 counter$count = 19288;
	#10 counter$count = 19289;
	#10 counter$count = 19290;
	#10 counter$count = 19291;
	#10 counter$count = 19292;
	#10 counter$count = 19293;
	#10 counter$count = 19294;
	#10 counter$count = 19295;
	#10 counter$count = 19296;
	#10 counter$count = 19297;
	#10 counter$count = 19298;
	#10 counter$count = 19299;
	#10 counter$count = 19300;
	#10 counter$count = 19301;
	#10 counter$count = 19302;
	#10 counter$count = 19303;
	#10 counter$count = 19304;
	#10 counter$count = 19305;
	#10 counter$count = 19306;
	#10 counter$count = 19307;
	#10 counter$count = 19308;
	#10 counter$count = 19309;
	#10 counter$count = 19310;
	#10 counter$count = 19311;
	#10 counter$count = 19312;
	#10 counter$count = 19313;
	#10 counter$count = 19314;
	#10 counter$count = 19315;
	#10 counter$count = 19316;
	#10 counter$count = 19317;
	#10 counter$count = 19318;
	#10 counter$count = 19319;
	#10 counter$count = 19320;
	#10 counter$count = 19321;
	#10 counter$count = 19322;
	#10 counter$count = 19323;
	#10 counter$count = 19324;
	#10 counter$count = 19325;
	#10 counter$count = 19326;
	#10 counter$count = 19327;
	#10 counter$count = 19328;
	#10 counter$count = 19329;
	#10 counter$count = 19330;
	#10 counter$count = 19331;
	#10 counter$count = 19332;
	#10 counter$count = 19333;
	#10 counter$count = 19334;
	#10 counter$count = 19335;
	#10 counter$count = 19336;
	#10 counter$count = 19337;
	#10 counter$count = 19338;
	#10 counter$count = 19339;
	#10 counter$count = 19340;
	#10 counter$count = 19341;
	#10 counter$count = 19342;
	#10 counter$count = 19343;
	#10 counter$count = 19344;
	#10 counter$count = 19345;
	#10 counter$count = 19346;
	#10 counter$count = 19347;
	#10 counter$count = 19348;
	#10 counter$count = 19349;
	#10 counter$count = 19350;
	#10 counter$count = 19351;
	#10 counter$count = 19352;
	#10 counter$count = 19353;
	#10 counter$count = 19354;
	#10 counter$count = 19355;
	#10 counter$count = 19356;
	#10 counter$count = 19357;
	#10 counter$count = 19358;
	#10 counter$count = 19359;
	#10 counter$count = 19360;
	#10 counter$count = 19361;
	#10 counter$count = 19362;
	#10 counter$count = 19363;
	#10 counter$count = 19364;
	#10 counter$count = 19365;
	#10 counter$count = 19366;
	#10 counter$count = 19367;
	#10 counter$count = 19368;
	#10 counter$count = 19369;
	#10 counter$count = 19370;
	#10 counter$count = 19371;
	#10 counter$count = 19372;
	#10 counter$count = 19373;
	#10 counter$count = 19374;
	#10 counter$count = 19375;
	#10 counter$count = 19376;
	#10 counter$count = 19377;
	#10 counter$count = 19378;
	#10 counter$count = 19379;
	#10 counter$count = 19380;
	#10 counter$count = 19381;
	#10 counter$count = 19382;
	#10 counter$count = 19383;
	#10 counter$count = 19384;
	#10 counter$count = 19385;
	#10 counter$count = 19386;
	#10 counter$count = 19387;
	#10 counter$count = 19388;
	#10 counter$count = 19389;
	#10 counter$count = 19390;
	#10 counter$count = 19391;
	#10 counter$count = 19392;
	#10 counter$count = 19393;
	#10 counter$count = 19394;
	#10 counter$count = 19395;
	#10 counter$count = 19396;
	#10 counter$count = 19397;
	#10 counter$count = 19398;
	#10 counter$count = 19399;
	#10 counter$count = 19400;
	#10 counter$count = 19401;
	#10 counter$count = 19402;
	#10 counter$count = 19403;
	#10 counter$count = 19404;
	#10 counter$count = 19405;
	#10 counter$count = 19406;
	#10 counter$count = 19407;
	#10 counter$count = 19408;
	#10 counter$count = 19409;
	#10 counter$count = 19410;
	#10 counter$count = 19411;
	#10 counter$count = 19412;
	#10 counter$count = 19413;
	#10 counter$count = 19414;
	#10 counter$count = 19415;
	#10 counter$count = 19416;
	#10 counter$count = 19417;
	#10 counter$count = 19418;
	#10 counter$count = 19419;
	#10 counter$count = 19420;
	#10 counter$count = 19421;
	#10 counter$count = 19422;
	#10 counter$count = 19423;
	#10 counter$count = 19424;
	#10 counter$count = 19425;
	#10 counter$count = 19426;
	#10 counter$count = 19427;
	#10 counter$count = 19428;
	#10 counter$count = 19429;
	#10 counter$count = 19430;
	#10 counter$count = 19431;
	#10 counter$count = 19432;
	#10 counter$count = 19433;
	#10 counter$count = 19434;
	#10 counter$count = 19435;
	#10 counter$count = 19436;
	#10 counter$count = 19437;
	#10 counter$count = 19438;
	#10 counter$count = 19439;
	#10 counter$count = 19440;
	#10 counter$count = 19441;
	#10 counter$count = 19442;
	#10 counter$count = 19443;
	#10 counter$count = 19444;
	#10 counter$count = 19445;
	#10 counter$count = 19446;
	#10 counter$count = 19447;
	#10 counter$count = 19448;
	#10 counter$count = 19449;
	#10 counter$count = 19450;
	#10 counter$count = 19451;
	#10 counter$count = 19452;
	#10 counter$count = 19453;
	#10 counter$count = 19454;
	#10 counter$count = 19455;
	#10 counter$count = 19456;
	#10 counter$count = 19457;
	#10 counter$count = 19458;
	#10 counter$count = 19459;
	#10 counter$count = 19460;
	#10 counter$count = 19461;
	#10 counter$count = 19462;
	#10 counter$count = 19463;
	#10 counter$count = 19464;
	#10 counter$count = 19465;
	#10 counter$count = 19466;
	#10 counter$count = 19467;
	#10 counter$count = 19468;
	#10 counter$count = 19469;
	#10 counter$count = 19470;
	#10 counter$count = 19471;
	#10 counter$count = 19472;
	#10 counter$count = 19473;
	#10 counter$count = 19474;
	#10 counter$count = 19475;
	#10 counter$count = 19476;
	#10 counter$count = 19477;
	#10 counter$count = 19478;
	#10 counter$count = 19479;
	#10 counter$count = 19480;
	#10 counter$count = 19481;
	#10 counter$count = 19482;
	#10 counter$count = 19483;
	#10 counter$count = 19484;
	#10 counter$count = 19485;
	#10 counter$count = 19486;
	#10 counter$count = 19487;
	#10 counter$count = 19488;
	#10 counter$count = 19489;
	#10 counter$count = 19490;
	#10 counter$count = 19491;
	#10 counter$count = 19492;
	#10 counter$count = 19493;
	#10 counter$count = 19494;
	#10 counter$count = 19495;
	#10 counter$count = 19496;
	#10 counter$count = 19497;
	#10 counter$count = 19498;
	#10 counter$count = 19499;
	#10 counter$count = 19500;
	#10 counter$count = 19501;
	#10 counter$count = 19502;
	#10 counter$count = 19503;
	#10 counter$count = 19504;
	#10 counter$count = 19505;
	#10 counter$count = 19506;
	#10 counter$count = 19507;
	#10 counter$count = 19508;
	#10 counter$count = 19509;
	#10 counter$count = 19510;
	#10 counter$count = 19511;
	#10 counter$count = 19512;
	#10 counter$count = 19513;
	#10 counter$count = 19514;
	#10 counter$count = 19515;
	#10 counter$count = 19516;
	#10 counter$count = 19517;
	#10 counter$count = 19518;
	#10 counter$count = 19519;
	#10 counter$count = 19520;
	#10 counter$count = 19521;
	#10 counter$count = 19522;
	#10 counter$count = 19523;
	#10 counter$count = 19524;
	#10 counter$count = 19525;
	#10 counter$count = 19526;
	#10 counter$count = 19527;
	#10 counter$count = 19528;
	#10 counter$count = 19529;
	#10 counter$count = 19530;
	#10 counter$count = 19531;
	#10 counter$count = 19532;
	#10 counter$count = 19533;
	#10 counter$count = 19534;
	#10 counter$count = 19535;
	#10 counter$count = 19536;
	#10 counter$count = 19537;
	#10 counter$count = 19538;
	#10 counter$count = 19539;
	#10 counter$count = 19540;
	#10 counter$count = 19541;
	#10 counter$count = 19542;
	#10 counter$count = 19543;
	#10 counter$count = 19544;
	#10 counter$count = 19545;
	#10 counter$count = 19546;
	#10 counter$count = 19547;
	#10 counter$count = 19548;
	#10 counter$count = 19549;
	#10 counter$count = 19550;
	#10 counter$count = 19551;
	#10 counter$count = 19552;
	#10 counter$count = 19553;
	#10 counter$count = 19554;
	#10 counter$count = 19555;
	#10 counter$count = 19556;
	#10 counter$count = 19557;
	#10 counter$count = 19558;
	#10 counter$count = 19559;
	#10 counter$count = 19560;
	#10 counter$count = 19561;
	#10 counter$count = 19562;
	#10 counter$count = 19563;
	#10 counter$count = 19564;
	#10 counter$count = 19565;
	#10 counter$count = 19566;
	#10 counter$count = 19567;
	#10 counter$count = 19568;
	#10 counter$count = 19569;
	#10 counter$count = 19570;
	#10 counter$count = 19571;
	#10 counter$count = 19572;
	#10 counter$count = 19573;
	#10 counter$count = 19574;
	#10 counter$count = 19575;
	#10 counter$count = 19576;
	#10 counter$count = 19577;
	#10 counter$count = 19578;
	#10 counter$count = 19579;
	#10 counter$count = 19580;
	#10 counter$count = 19581;
	#10 counter$count = 19582;
	#10 counter$count = 19583;
	#10 counter$count = 19584;
	#10 counter$count = 19585;
	#10 counter$count = 19586;
	#10 counter$count = 19587;
	#10 counter$count = 19588;
	#10 counter$count = 19589;
	#10 counter$count = 19590;
	#10 counter$count = 19591;
	#10 counter$count = 19592;
	#10 counter$count = 19593;
	#10 counter$count = 19594;
	#10 counter$count = 19595;
	#10 counter$count = 19596;
	#10 counter$count = 19597;
	#10 counter$count = 19598;
	#10 counter$count = 19599;
	#10 counter$count = 19600;
	#10 counter$count = 19601;
	#10 counter$count = 19602;
	#10 counter$count = 19603;
	#10 counter$count = 19604;
	#10 counter$count = 19605;
	#10 counter$count = 19606;
	#10 counter$count = 19607;
	#10 counter$count = 19608;
	#10 counter$count = 19609;
	#10 counter$count = 19610;
	#10 counter$count = 19611;
	#10 counter$count = 19612;
	#10 counter$count = 19613;
	#10 counter$count = 19614;
	#10 counter$count = 19615;
	#10 counter$count = 19616;
	#10 counter$count = 19617;
	#10 counter$count = 19618;
	#10 counter$count = 19619;
	#10 counter$count = 19620;
	#10 counter$count = 19621;
	#10 counter$count = 19622;
	#10 counter$count = 19623;
	#10 counter$count = 19624;
	#10 counter$count = 19625;
	#10 counter$count = 19626;
	#10 counter$count = 19627;
	#10 counter$count = 19628;
	#10 counter$count = 19629;
	#10 counter$count = 19630;
	#10 counter$count = 19631;
	#10 counter$count = 19632;
	#10 counter$count = 19633;
	#10 counter$count = 19634;
	#10 counter$count = 19635;
	#10 counter$count = 19636;
	#10 counter$count = 19637;
	#10 counter$count = 19638;
	#10 counter$count = 19639;
	#10 counter$count = 19640;
	#10 counter$count = 19641;
	#10 counter$count = 19642;
	#10 counter$count = 19643;
	#10 counter$count = 19644;
	#10 counter$count = 19645;
	#10 counter$count = 19646;
	#10 counter$count = 19647;
	#10 counter$count = 19648;
	#10 counter$count = 19649;
	#10 counter$count = 19650;
	#10 counter$count = 19651;
	#10 counter$count = 19652;
	#10 counter$count = 19653;
	#10 counter$count = 19654;
	#10 counter$count = 19655;
	#10 counter$count = 19656;
	#10 counter$count = 19657;
	#10 counter$count = 19658;
	#10 counter$count = 19659;
	#10 counter$count = 19660;
	#10 counter$count = 19661;
	#10 counter$count = 19662;
	#10 counter$count = 19663;
	#10 counter$count = 19664;
	#10 counter$count = 19665;
	#10 counter$count = 19666;
	#10 counter$count = 19667;
	#10 counter$count = 19668;
	#10 counter$count = 19669;
	#10 counter$count = 19670;
	#10 counter$count = 19671;
	#10 counter$count = 19672;
	#10 counter$count = 19673;
	#10 counter$count = 19674;
	#10 counter$count = 19675;
	#10 counter$count = 19676;
	#10 counter$count = 19677;
	#10 counter$count = 19678;
	#10 counter$count = 19679;
	#10 counter$count = 19680;
	#10 counter$count = 19681;
	#10 counter$count = 19682;
	#10 counter$count = 19683;
	#10 counter$count = 19684;
	#10 counter$count = 19685;
	#10 counter$count = 19686;
	#10 counter$count = 19687;
	#10 counter$count = 19688;
	#10 counter$count = 19689;
	#10 counter$count = 19690;
	#10 counter$count = 19691;
	#10 counter$count = 19692;
	#10 counter$count = 19693;
	#10 counter$count = 19694;
	#10 counter$count = 19695;
	#10 counter$count = 19696;
	#10 counter$count = 19697;
	#10 counter$count = 19698;
	#10 counter$count = 19699;
	#10 counter$count = 19700;
	#10 counter$count = 19701;
	#10 counter$count = 19702;
	#10 counter$count = 19703;
	#10 counter$count = 19704;
	#10 counter$count = 19705;
	#10 counter$count = 19706;
	#10 counter$count = 19707;
	#10 counter$count = 19708;
	#10 counter$count = 19709;
	#10 counter$count = 19710;
	#10 counter$count = 19711;
	#10 counter$count = 19712;
	#10 counter$count = 19713;
	#10 counter$count = 19714;
	#10 counter$count = 19715;
	#10 counter$count = 19716;
	#10 counter$count = 19717;
	#10 counter$count = 19718;
	#10 counter$count = 19719;
	#10 counter$count = 19720;
	#10 counter$count = 19721;
	#10 counter$count = 19722;
	#10 counter$count = 19723;
	#10 counter$count = 19724;
	#10 counter$count = 19725;
	#10 counter$count = 19726;
	#10 counter$count = 19727;
	#10 counter$count = 19728;
	#10 counter$count = 19729;
	#10 counter$count = 19730;
	#10 counter$count = 19731;
	#10 counter$count = 19732;
	#10 counter$count = 19733;
	#10 counter$count = 19734;
	#10 counter$count = 19735;
	#10 counter$count = 19736;
	#10 counter$count = 19737;
	#10 counter$count = 19738;
	#10 counter$count = 19739;
	#10 counter$count = 19740;
	#10 counter$count = 19741;
	#10 counter$count = 19742;
	#10 counter$count = 19743;
	#10 counter$count = 19744;
	#10 counter$count = 19745;
	#10 counter$count = 19746;
	#10 counter$count = 19747;
	#10 counter$count = 19748;
	#10 counter$count = 19749;
	#10 counter$count = 19750;
	#10 counter$count = 19751;
	#10 counter$count = 19752;
	#10 counter$count = 19753;
	#10 counter$count = 19754;
	#10 counter$count = 19755;
	#10 counter$count = 19756;
	#10 counter$count = 19757;
	#10 counter$count = 19758;
	#10 counter$count = 19759;
	#10 counter$count = 19760;
	#10 counter$count = 19761;
	#10 counter$count = 19762;
	#10 counter$count = 19763;
	#10 counter$count = 19764;
	#10 counter$count = 19765;
	#10 counter$count = 19766;
	#10 counter$count = 19767;
	#10 counter$count = 19768;
	#10 counter$count = 19769;
	#10 counter$count = 19770;
	#10 counter$count = 19771;
	#10 counter$count = 19772;
	#10 counter$count = 19773;
	#10 counter$count = 19774;
	#10 counter$count = 19775;
	#10 counter$count = 19776;
	#10 counter$count = 19777;
	#10 counter$count = 19778;
	#10 counter$count = 19779;
	#10 counter$count = 19780;
	#10 counter$count = 19781;
	#10 counter$count = 19782;
	#10 counter$count = 19783;
	#10 counter$count = 19784;
	#10 counter$count = 19785;
	#10 counter$count = 19786;
	#10 counter$count = 19787;
	#10 counter$count = 19788;
	#10 counter$count = 19789;
	#10 counter$count = 19790;
	#10 counter$count = 19791;
	#10 counter$count = 19792;
	#10 counter$count = 19793;
	#10 counter$count = 19794;
	#10 counter$count = 19795;
	#10 counter$count = 19796;
	#10 counter$count = 19797;
	#10 counter$count = 19798;
	#10 counter$count = 19799;
	#10 counter$count = 19800;
	#10 counter$count = 19801;
	#10 counter$count = 19802;
	#10 counter$count = 19803;
	#10 counter$count = 19804;
	#10 counter$count = 19805;
	#10 counter$count = 19806;
	#10 counter$count = 19807;
	#10 counter$count = 19808;
	#10 counter$count = 19809;
	#10 counter$count = 19810;
	#10 counter$count = 19811;
	#10 counter$count = 19812;
	#10 counter$count = 19813;
	#10 counter$count = 19814;
	#10 counter$count = 19815;
	#10 counter$count = 19816;
	#10 counter$count = 19817;
	#10 counter$count = 19818;
	#10 counter$count = 19819;
	#10 counter$count = 19820;
	#10 counter$count = 19821;
	#10 counter$count = 19822;
	#10 counter$count = 19823;
	#10 counter$count = 19824;
	#10 counter$count = 19825;
	#10 counter$count = 19826;
	#10 counter$count = 19827;
	#10 counter$count = 19828;
	#10 counter$count = 19829;
	#10 counter$count = 19830;
	#10 counter$count = 19831;
	#10 counter$count = 19832;
	#10 counter$count = 19833;
	#10 counter$count = 19834;
	#10 counter$count = 19835;
	#10 counter$count = 19836;
	#10 counter$count = 19837;
	#10 counter$count = 19838;
	#10 counter$count = 19839;
	#10 counter$count = 19840;
	#10 counter$count = 19841;
	#10 counter$count = 19842;
	#10 counter$count = 19843;
	#10 counter$count = 19844;
	#10 counter$count = 19845;
	#10 counter$count = 19846;
	#10 counter$count = 19847;
	#10 counter$count = 19848;
	#10 counter$count = 19849;
	#10 counter$count = 19850;
	#10 counter$count = 19851;
	#10 counter$count = 19852;
	#10 counter$count = 19853;
	#10 counter$count = 19854;
	#10 counter$count = 19855;
	#10 counter$count = 19856;
	#10 counter$count = 19857;
	#10 counter$count = 19858;
	#10 counter$count = 19859;
	#10 counter$count = 19860;
	#10 counter$count = 19861;
	#10 counter$count = 19862;
	#10 counter$count = 19863;
	#10 counter$count = 19864;
	#10 counter$count = 19865;
	#10 counter$count = 19866;
	#10 counter$count = 19867;
	#10 counter$count = 19868;
	#10 counter$count = 19869;
	#10 counter$count = 19870;
	#10 counter$count = 19871;
	#10 counter$count = 19872;
	#10 counter$count = 19873;
	#10 counter$count = 19874;
	#10 counter$count = 19875;
	#10 counter$count = 19876;
	#10 counter$count = 19877;
	#10 counter$count = 19878;
	#10 counter$count = 19879;
	#10 counter$count = 19880;
	#10 counter$count = 19881;
	#10 counter$count = 19882;
	#10 counter$count = 19883;
	#10 counter$count = 19884;
	#10 counter$count = 19885;
	#10 counter$count = 19886;
	#10 counter$count = 19887;
	#10 counter$count = 19888;
	#10 counter$count = 19889;
	#10 counter$count = 19890;
	#10 counter$count = 19891;
	#10 counter$count = 19892;
	#10 counter$count = 19893;
	#10 counter$count = 19894;
	#10 counter$count = 19895;
	#10 counter$count = 19896;
	#10 counter$count = 19897;
	#10 counter$count = 19898;
	#10 counter$count = 19899;
	#10 counter$count = 19900;
	#10 counter$count = 19901;
	#10 counter$count = 19902;
	#10 counter$count = 19903;
	#10 counter$count = 19904;
	#10 counter$count = 19905;
	#10 counter$count = 19906;
	#10 counter$count = 19907;
	#10 counter$count = 19908;
	#10 counter$count = 19909;
	#10 counter$count = 19910;
	#10 counter$count = 19911;
	#10 counter$count = 19912;
	#10 counter$count = 19913;
	#10 counter$count = 19914;
	#10 counter$count = 19915;
	#10 counter$count = 19916;
	#10 counter$count = 19917;
	#10 counter$count = 19918;
	#10 counter$count = 19919;
	#10 counter$count = 19920;
	#10 counter$count = 19921;
	#10 counter$count = 19922;
	#10 counter$count = 19923;
	#10 counter$count = 19924;
	#10 counter$count = 19925;
	#10 counter$count = 19926;
	#10 counter$count = 19927;
	#10 counter$count = 19928;
	#10 counter$count = 19929;
	#10 counter$count = 19930;
	#10 counter$count = 19931;
	#10 counter$count = 19932;
	#10 counter$count = 19933;
	#10 counter$count = 19934;
	#10 counter$count = 19935;
	#10 counter$count = 19936;
	#10 counter$count = 19937;
	#10 counter$count = 19938;
	#10 counter$count = 19939;
	#10 counter$count = 19940;
	#10 counter$count = 19941;
	#10 counter$count = 19942;
	#10 counter$count = 19943;
	#10 counter$count = 19944;
	#10 counter$count = 19945;
	#10 counter$count = 19946;
	#10 counter$count = 19947;
	#10 counter$count = 19948;
	#10 counter$count = 19949;
	#10 counter$count = 19950;
	#10 counter$count = 19951;
	#10 counter$count = 19952;
	#10 counter$count = 19953;
	#10 counter$count = 19954;
	#10 counter$count = 19955;
	#10 counter$count = 19956;
	#10 counter$count = 19957;
	#10 counter$count = 19958;
	#10 counter$count = 19959;
	#10 counter$count = 19960;
	#10 counter$count = 19961;
	#10 counter$count = 19962;
	#10 counter$count = 19963;
	#10 counter$count = 19964;
	#10 counter$count = 19965;
	#10 counter$count = 19966;
	#10 counter$count = 19967;
	#10 counter$count = 19968;
	#10 counter$count = 19969;
	#10 counter$count = 19970;
	#10 counter$count = 19971;
	#10 counter$count = 19972;
	#10 counter$count = 19973;
	#10 counter$count = 19974;
	#10 counter$count = 19975;
	#10 counter$count = 19976;
	#10 counter$count = 19977;
	#10 counter$count = 19978;
	#10 counter$count = 19979;
	#10 counter$count = 19980;
	#10 counter$count = 19981;
	#10 counter$count = 19982;
	#10 counter$count = 19983;
	#10 counter$count = 19984;
	#10 counter$count = 19985;
	#10 counter$count = 19986;
	#10 counter$count = 19987;
	#10 counter$count = 19988;
	#10 counter$count = 19989;
	#10 counter$count = 19990;
	#10 counter$count = 19991;
	#10 counter$count = 19992;
	#10 counter$count = 19993;
	#10 counter$count = 19994;
	#10 counter$count = 19995;
	#10 counter$count = 19996;
	#10 counter$count = 19997;
	#10 counter$count = 19998;
	#10 counter$count = 19999;
	#10 counter$count = 20000;
	#10 counter$count = 20001;
	#10 counter$count = 20002;
	#10 counter$count = 20003;
	#10 counter$count = 20004;
	#10 counter$count = 20005;
	#10 counter$count = 20006;
	#10 counter$count = 20007;
	#10 counter$count = 20008;
	#10 counter$count = 20009;
	#10 counter$count = 20010;
	#10 counter$count = 20011;
	#10 counter$count = 20012;
	#10 counter$count = 20013;
	#10 counter$count = 20014;
	#10 counter$count = 20015;
	#10 counter$count = 20016;
	#10 counter$count = 20017;
	#10 counter$count = 20018;
	#10 counter$count = 20019;
	#10 counter$count = 20020;
	#10 counter$count = 20021;
	#10 counter$count = 20022;
	#10 counter$count = 20023;
	#10 counter$count = 20024;
	#10 counter$count = 20025;
	#10 counter$count = 20026;
	#10 counter$count = 20027;
	#10 counter$count = 20028;
	#10 counter$count = 20029;
	#10 counter$count = 20030;
	#10 counter$count = 20031;
	#10 counter$count = 20032;
	#10 counter$count = 20033;
	#10 counter$count = 20034;
	#10 counter$count = 20035;
	#10 counter$count = 20036;
	#10 counter$count = 20037;
	#10 counter$count = 20038;
	#10 counter$count = 20039;
	#10 counter$count = 20040;
	#10 counter$count = 20041;
	#10 counter$count = 20042;
	#10 counter$count = 20043;
	#10 counter$count = 20044;
	#10 counter$count = 20045;
	#10 counter$count = 20046;
	#10 counter$count = 20047;
	#10 counter$count = 20048;
	#10 counter$count = 20049;
	#10 counter$count = 20050;
	#10 counter$count = 20051;
	#10 counter$count = 20052;
	#10 counter$count = 20053;
	#10 counter$count = 20054;
	#10 counter$count = 20055;
	#10 counter$count = 20056;
	#10 counter$count = 20057;
	#10 counter$count = 20058;
	#10 counter$count = 20059;
	#10 counter$count = 20060;
	#10 counter$count = 20061;
	#10 counter$count = 20062;
	#10 counter$count = 20063;
	#10 counter$count = 20064;
	#10 counter$count = 20065;
	#10 counter$count = 20066;
	#10 counter$count = 20067;
	#10 counter$count = 20068;
	#10 counter$count = 20069;
	#10 counter$count = 20070;
	#10 counter$count = 20071;
	#10 counter$count = 20072;
	#10 counter$count = 20073;
	#10 counter$count = 20074;
	#10 counter$count = 20075;
	#10 counter$count = 20076;
	#10 counter$count = 20077;
	#10 counter$count = 20078;
	#10 counter$count = 20079;
	#10 counter$count = 20080;
	#10 counter$count = 20081;
	#10 counter$count = 20082;
	#10 counter$count = 20083;
	#10 counter$count = 20084;
	#10 counter$count = 20085;
	#10 counter$count = 20086;
	#10 counter$count = 20087;
	#10 counter$count = 20088;
	#10 counter$count = 20089;
	#10 counter$count = 20090;
	#10 counter$count = 20091;
	#10 counter$count = 20092;
	#10 counter$count = 20093;
	#10 counter$count = 20094;
	#10 counter$count = 20095;
	#10 counter$count = 20096;
	#10 counter$count = 20097;
	#10 counter$count = 20098;
	#10 counter$count = 20099;
	#10 counter$count = 20100;
	#10 counter$count = 20101;
	#10 counter$count = 20102;
	#10 counter$count = 20103;
	#10 counter$count = 20104;
	#10 counter$count = 20105;
	#10 counter$count = 20106;
	#10 counter$count = 20107;
	#10 counter$count = 20108;
	#10 counter$count = 20109;
	#10 counter$count = 20110;
	#10 counter$count = 20111;
	#10 counter$count = 20112;
	#10 counter$count = 20113;
	#10 counter$count = 20114;
	#10 counter$count = 20115;
	#10 counter$count = 20116;
	#10 counter$count = 20117;
	#10 counter$count = 20118;
	#10 counter$count = 20119;
	#10 counter$count = 20120;
	#10 counter$count = 20121;
	#10 counter$count = 20122;
	#10 counter$count = 20123;
	#10 counter$count = 20124;
	#10 counter$count = 20125;
	#10 counter$count = 20126;
	#10 counter$count = 20127;
	#10 counter$count = 20128;
	#10 counter$count = 20129;
	#10 counter$count = 20130;
	#10 counter$count = 20131;
	#10 counter$count = 20132;
	#10 counter$count = 20133;
	#10 counter$count = 20134;
	#10 counter$count = 20135;
	#10 counter$count = 20136;
	#10 counter$count = 20137;
	#10 counter$count = 20138;
	#10 counter$count = 20139;
	#10 counter$count = 20140;
	#10 counter$count = 20141;
	#10 counter$count = 20142;
	#10 counter$count = 20143;
	#10 counter$count = 20144;
	#10 counter$count = 20145;
	#10 counter$count = 20146;
	#10 counter$count = 20147;
	#10 counter$count = 20148;
	#10 counter$count = 20149;
	#10 counter$count = 20150;
	#10 counter$count = 20151;
	#10 counter$count = 20152;
	#10 counter$count = 20153;
	#10 counter$count = 20154;
	#10 counter$count = 20155;
	#10 counter$count = 20156;
	#10 counter$count = 20157;
	#10 counter$count = 20158;
	#10 counter$count = 20159;
	#10 counter$count = 20160;
	#10 counter$count = 20161;
	#10 counter$count = 20162;
	#10 counter$count = 20163;
	#10 counter$count = 20164;
	#10 counter$count = 20165;
	#10 counter$count = 20166;
	#10 counter$count = 20167;
	#10 counter$count = 20168;
	#10 counter$count = 20169;
	#10 counter$count = 20170;
	#10 counter$count = 20171;
	#10 counter$count = 20172;
	#10 counter$count = 20173;
	#10 counter$count = 20174;
	#10 counter$count = 20175;
	#10 counter$count = 20176;
	#10 counter$count = 20177;
	#10 counter$count = 20178;
	#10 counter$count = 20179;
	#10 counter$count = 20180;
	#10 counter$count = 20181;
	#10 counter$count = 20182;
	#10 counter$count = 20183;
	#10 counter$count = 20184;
	#10 counter$count = 20185;
	#10 counter$count = 20186;
	#10 counter$count = 20187;
	#10 counter$count = 20188;
	#10 counter$count = 20189;
	#10 counter$count = 20190;
	#10 counter$count = 20191;
	#10 counter$count = 20192;
	#10 counter$count = 20193;
	#10 counter$count = 20194;
	#10 counter$count = 20195;
	#10 counter$count = 20196;
	#10 counter$count = 20197;
	#10 counter$count = 20198;
	#10 counter$count = 20199;
	#10 counter$count = 20200;
	#10 counter$count = 20201;
	#10 counter$count = 20202;
	#10 counter$count = 20203;
	#10 counter$count = 20204;
	#10 counter$count = 20205;
	#10 counter$count = 20206;
	#10 counter$count = 20207;
	#10 counter$count = 20208;
	#10 counter$count = 20209;
	#10 counter$count = 20210;
	#10 counter$count = 20211;
	#10 counter$count = 20212;
	#10 counter$count = 20213;
	#10 counter$count = 20214;
	#10 counter$count = 20215;
	#10 counter$count = 20216;
	#10 counter$count = 20217;
	#10 counter$count = 20218;
	#10 counter$count = 20219;
	#10 counter$count = 20220;
	#10 counter$count = 20221;
	#10 counter$count = 20222;
	#10 counter$count = 20223;
	#10 counter$count = 20224;
	#10 counter$count = 20225;
	#10 counter$count = 20226;
	#10 counter$count = 20227;
	#10 counter$count = 20228;
	#10 counter$count = 20229;
	#10 counter$count = 20230;
	#10 counter$count = 20231;
	#10 counter$count = 20232;
	#10 counter$count = 20233;
	#10 counter$count = 20234;
	#10 counter$count = 20235;
	#10 counter$count = 20236;
	#10 counter$count = 20237;
	#10 counter$count = 20238;
	#10 counter$count = 20239;
	#10 counter$count = 20240;
	#10 counter$count = 20241;
	#10 counter$count = 20242;
	#10 counter$count = 20243;
	#10 counter$count = 20244;
	#10 counter$count = 20245;
	#10 counter$count = 20246;
	#10 counter$count = 20247;
	#10 counter$count = 20248;
	#10 counter$count = 20249;
	#10 counter$count = 20250;
	#10 counter$count = 20251;
	#10 counter$count = 20252;
	#10 counter$count = 20253;
	#10 counter$count = 20254;
	#10 counter$count = 20255;
	#10 counter$count = 20256;
	#10 counter$count = 20257;
	#10 counter$count = 20258;
	#10 counter$count = 20259;
	#10 counter$count = 20260;
	#10 counter$count = 20261;
	#10 counter$count = 20262;
	#10 counter$count = 20263;
	#10 counter$count = 20264;
	#10 counter$count = 20265;
	#10 counter$count = 20266;
	#10 counter$count = 20267;
	#10 counter$count = 20268;
	#10 counter$count = 20269;
	#10 counter$count = 20270;
	#10 counter$count = 20271;
	#10 counter$count = 20272;
	#10 counter$count = 20273;
	#10 counter$count = 20274;
	#10 counter$count = 20275;
	#10 counter$count = 20276;
	#10 counter$count = 20277;
	#10 counter$count = 20278;
	#10 counter$count = 20279;
	#10 counter$count = 20280;
	#10 counter$count = 20281;
	#10 counter$count = 20282;
	#10 counter$count = 20283;
	#10 counter$count = 20284;
	#10 counter$count = 20285;
	#10 counter$count = 20286;
	#10 counter$count = 20287;
	#10 counter$count = 20288;
	#10 counter$count = 20289;
	#10 counter$count = 20290;
	#10 counter$count = 20291;
	#10 counter$count = 20292;
	#10 counter$count = 20293;
	#10 counter$count = 20294;
	#10 counter$count = 20295;
	#10 counter$count = 20296;
	#10 counter$count = 20297;
	#10 counter$count = 20298;
	#10 counter$count = 20299;
	#10 counter$count = 20300;
	#10 counter$count = 20301;
	#10 counter$count = 20302;
	#10 counter$count = 20303;
	#10 counter$count = 20304;
	#10 counter$count = 20305;
	#10 counter$count = 20306;
	#10 counter$count = 20307;
	#10 counter$count = 20308;
	#10 counter$count = 20309;
	#10 counter$count = 20310;
	#10 counter$count = 20311;
	#10 counter$count = 20312;
	#10 counter$count = 20313;
	#10 counter$count = 20314;
	#10 counter$count = 20315;
	#10 counter$count = 20316;
	#10 counter$count = 20317;
	#10 counter$count = 20318;
	#10 counter$count = 20319;
	#10 counter$count = 20320;
	#10 counter$count = 20321;
	#10 counter$count = 20322;
	#10 counter$count = 20323;
	#10 counter$count = 20324;
	#10 counter$count = 20325;
	#10 counter$count = 20326;
	#10 counter$count = 20327;
	#10 counter$count = 20328;
	#10 counter$count = 20329;
	#10 counter$count = 20330;
	#10 counter$count = 20331;
	#10 counter$count = 20332;
	#10 counter$count = 20333;
	#10 counter$count = 20334;
	#10 counter$count = 20335;
	#10 counter$count = 20336;
	#10 counter$count = 20337;
	#10 counter$count = 20338;
	#10 counter$count = 20339;
	#10 counter$count = 20340;
	#10 counter$count = 20341;
	#10 counter$count = 20342;
	#10 counter$count = 20343;
	#10 counter$count = 20344;
	#10 counter$count = 20345;
	#10 counter$count = 20346;
	#10 counter$count = 20347;
	#10 counter$count = 20348;
	#10 counter$count = 20349;
	#10 counter$count = 20350;
	#10 counter$count = 20351;
	#10 counter$count = 20352;
	#10 counter$count = 20353;
	#10 counter$count = 20354;
	#10 counter$count = 20355;
	#10 counter$count = 20356;
	#10 counter$count = 20357;
	#10 counter$count = 20358;
	#10 counter$count = 20359;
	#10 counter$count = 20360;
	#10 counter$count = 20361;
	#10 counter$count = 20362;
	#10 counter$count = 20363;
	#10 counter$count = 20364;
	#10 counter$count = 20365;
	#10 counter$count = 20366;
	#10 counter$count = 20367;
	#10 counter$count = 20368;
	#10 counter$count = 20369;
	#10 counter$count = 20370;
	#10 counter$count = 20371;
	#10 counter$count = 20372;
	#10 counter$count = 20373;
	#10 counter$count = 20374;
	#10 counter$count = 20375;
	#10 counter$count = 20376;
	#10 counter$count = 20377;
	#10 counter$count = 20378;
	#10 counter$count = 20379;
	#10 counter$count = 20380;
	#10 counter$count = 20381;
	#10 counter$count = 20382;
	#10 counter$count = 20383;
	#10 counter$count = 20384;
	#10 counter$count = 20385;
	#10 counter$count = 20386;
	#10 counter$count = 20387;
	#10 counter$count = 20388;
	#10 counter$count = 20389;
	#10 counter$count = 20390;
	#10 counter$count = 20391;
	#10 counter$count = 20392;
	#10 counter$count = 20393;
	#10 counter$count = 20394;
	#10 counter$count = 20395;
	#10 counter$count = 20396;
	#10 counter$count = 20397;
	#10 counter$count = 20398;
	#10 counter$count = 20399;
	#10 counter$count = 20400;
	#10 counter$count = 20401;
	#10 counter$count = 20402;
	#10 counter$count = 20403;
	#10 counter$count = 20404;
	#10 counter$count = 20405;
	#10 counter$count = 20406;
	#10 counter$count = 20407;
	#10 counter$count = 20408;
	#10 counter$count = 20409;
	#10 counter$count = 20410;
	#10 counter$count = 20411;
	#10 counter$count = 20412;
	#10 counter$count = 20413;
	#10 counter$count = 20414;
	#10 counter$count = 20415;
	#10 counter$count = 20416;
	#10 counter$count = 20417;
	#10 counter$count = 20418;
	#10 counter$count = 20419;
	#10 counter$count = 20420;
	#10 counter$count = 20421;
	#10 counter$count = 20422;
	#10 counter$count = 20423;
	#10 counter$count = 20424;
	#10 counter$count = 20425;
	#10 counter$count = 20426;
	#10 counter$count = 20427;
	#10 counter$count = 20428;
	#10 counter$count = 20429;
	#10 counter$count = 20430;
	#10 counter$count = 20431;
	#10 counter$count = 20432;
	#10 counter$count = 20433;
	#10 counter$count = 20434;
	#10 counter$count = 20435;
	#10 counter$count = 20436;
	#10 counter$count = 20437;
	#10 counter$count = 20438;
	#10 counter$count = 20439;
	#10 counter$count = 20440;
	#10 counter$count = 20441;
	#10 counter$count = 20442;
	#10 counter$count = 20443;
	#10 counter$count = 20444;
	#10 counter$count = 20445;
	#10 counter$count = 20446;
	#10 counter$count = 20447;
	#10 counter$count = 20448;
	#10 counter$count = 20449;
	#10 counter$count = 20450;
	#10 counter$count = 20451;
	#10 counter$count = 20452;
	#10 counter$count = 20453;
	#10 counter$count = 20454;
	#10 counter$count = 20455;
	#10 counter$count = 20456;
	#10 counter$count = 20457;
	#10 counter$count = 20458;
	#10 counter$count = 20459;
	#10 counter$count = 20460;
	#10 counter$count = 20461;
	#10 counter$count = 20462;
	#10 counter$count = 20463;
	#10 counter$count = 20464;
	#10 counter$count = 20465;
	#10 counter$count = 20466;
	#10 counter$count = 20467;
	#10 counter$count = 20468;
	#10 counter$count = 20469;
	#10 counter$count = 20470;
	#10 counter$count = 20471;
	#10 counter$count = 20472;
	#10 counter$count = 20473;
	#10 counter$count = 20474;
	#10 counter$count = 20475;
	#10 counter$count = 20476;
	#10 counter$count = 20477;
	#10 counter$count = 20478;
	#10 counter$count = 20479;
	#10 counter$count = 20480;
	#10 counter$count = 20481;
	#10 counter$count = 20482;
	#10 counter$count = 20483;
	#10 counter$count = 20484;
	#10 counter$count = 20485;
	#10 counter$count = 20486;
	#10 counter$count = 20487;
	#10 counter$count = 20488;
	#10 counter$count = 20489;
	#10 counter$count = 20490;
	#10 counter$count = 20491;
	#10 counter$count = 20492;
	#10 counter$count = 20493;
	#10 counter$count = 20494;
	#10 counter$count = 20495;
	#10 counter$count = 20496;
	#10 counter$count = 20497;
	#10 counter$count = 20498;
	#10 counter$count = 20499;
	#10 counter$count = 20500;
	#10 counter$count = 20501;
	#10 counter$count = 20502;
	#10 counter$count = 20503;
	#10 counter$count = 20504;
	#10 counter$count = 20505;
	#10 counter$count = 20506;
	#10 counter$count = 20507;
	#10 counter$count = 20508;
	#10 counter$count = 20509;
	#10 counter$count = 20510;
	#10 counter$count = 20511;
	#10 counter$count = 20512;
	#10 counter$count = 20513;
	#10 counter$count = 20514;
	#10 counter$count = 20515;
	#10 counter$count = 20516;
	#10 counter$count = 20517;
	#10 counter$count = 20518;
	#10 counter$count = 20519;
	#10 counter$count = 20520;
	#10 counter$count = 20521;
	#10 counter$count = 20522;
	#10 counter$count = 20523;
	#10 counter$count = 20524;
	#10 counter$count = 20525;
	#10 counter$count = 20526;
	#10 counter$count = 20527;
	#10 counter$count = 20528;
	#10 counter$count = 20529;
	#10 counter$count = 20530;
	#10 counter$count = 20531;
	#10 counter$count = 20532;
	#10 counter$count = 20533;
	#10 counter$count = 20534;
	#10 counter$count = 20535;
	#10 counter$count = 20536;
	#10 counter$count = 20537;
	#10 counter$count = 20538;
	#10 counter$count = 20539;
	#10 counter$count = 20540;
	#10 counter$count = 20541;
	#10 counter$count = 20542;
	#10 counter$count = 20543;
	#10 counter$count = 20544;
	#10 counter$count = 20545;
	#10 counter$count = 20546;
	#10 counter$count = 20547;
	#10 counter$count = 20548;
	#10 counter$count = 20549;
	#10 counter$count = 20550;
	#10 counter$count = 20551;
	#10 counter$count = 20552;
	#10 counter$count = 20553;
	#10 counter$count = 20554;
	#10 counter$count = 20555;
	#10 counter$count = 20556;
	#10 counter$count = 20557;
	#10 counter$count = 20558;
	#10 counter$count = 20559;
	#10 counter$count = 20560;
	#10 counter$count = 20561;
	#10 counter$count = 20562;
	#10 counter$count = 20563;
	#10 counter$count = 20564;
	#10 counter$count = 20565;
	#10 counter$count = 20566;
	#10 counter$count = 20567;
	#10 counter$count = 20568;
	#10 counter$count = 20569;
	#10 counter$count = 20570;
	#10 counter$count = 20571;
	#10 counter$count = 20572;
	#10 counter$count = 20573;
	#10 counter$count = 20574;
	#10 counter$count = 20575;
	#10 counter$count = 20576;
	#10 counter$count = 20577;
	#10 counter$count = 20578;
	#10 counter$count = 20579;
	#10 counter$count = 20580;
	#10 counter$count = 20581;
	#10 counter$count = 20582;
	#10 counter$count = 20583;
	#10 counter$count = 20584;
	#10 counter$count = 20585;
	#10 counter$count = 20586;
	#10 counter$count = 20587;
	#10 counter$count = 20588;
	#10 counter$count = 20589;
	#10 counter$count = 20590;
	#10 counter$count = 20591;
	#10 counter$count = 20592;
	#10 counter$count = 20593;
	#10 counter$count = 20594;
	#10 counter$count = 20595;
	#10 counter$count = 20596;
	#10 counter$count = 20597;
	#10 counter$count = 20598;
	#10 counter$count = 20599;
	#10 counter$count = 20600;
	#10 counter$count = 20601;
	#10 counter$count = 20602;
	#10 counter$count = 20603;
	#10 counter$count = 20604;
	#10 counter$count = 20605;
	#10 counter$count = 20606;
	#10 counter$count = 20607;
	#10 counter$count = 20608;
	#10 counter$count = 20609;
	#10 counter$count = 20610;
	#10 counter$count = 20611;
	#10 counter$count = 20612;
	#10 counter$count = 20613;
	#10 counter$count = 20614;
	#10 counter$count = 20615;
	#10 counter$count = 20616;
	#10 counter$count = 20617;
	#10 counter$count = 20618;
	#10 counter$count = 20619;
	#10 counter$count = 20620;
	#10 counter$count = 20621;
	#10 counter$count = 20622;
	#10 counter$count = 20623;
	#10 counter$count = 20624;
	#10 counter$count = 20625;
	#10 counter$count = 20626;
	#10 counter$count = 20627;
	#10 counter$count = 20628;
	#10 counter$count = 20629;
	#10 counter$count = 20630;
	#10 counter$count = 20631;
	#10 counter$count = 20632;
	#10 counter$count = 20633;
	#10 counter$count = 20634;
	#10 counter$count = 20635;
	#10 counter$count = 20636;
	#10 counter$count = 20637;
	#10 counter$count = 20638;
	#10 counter$count = 20639;
	#10 counter$count = 20640;
	#10 counter$count = 20641;
	#10 counter$count = 20642;
	#10 counter$count = 20643;
	#10 counter$count = 20644;
	#10 counter$count = 20645;
	#10 counter$count = 20646;
	#10 counter$count = 20647;
	#10 counter$count = 20648;
	#10 counter$count = 20649;
	#10 counter$count = 20650;
	#10 counter$count = 20651;
	#10 counter$count = 20652;
	#10 counter$count = 20653;
	#10 counter$count = 20654;
	#10 counter$count = 20655;
	#10 counter$count = 20656;
	#10 counter$count = 20657;
	#10 counter$count = 20658;
	#10 counter$count = 20659;
	#10 counter$count = 20660;
	#10 counter$count = 20661;
	#10 counter$count = 20662;
	#10 counter$count = 20663;
	#10 counter$count = 20664;
	#10 counter$count = 20665;
	#10 counter$count = 20666;
	#10 counter$count = 20667;
	#10 counter$count = 20668;
	#10 counter$count = 20669;
	#10 counter$count = 20670;
	#10 counter$count = 20671;
	#10 counter$count = 20672;
	#10 counter$count = 20673;
	#10 counter$count = 20674;
	#10 counter$count = 20675;
	#10 counter$count = 20676;
	#10 counter$count = 20677;
	#10 counter$count = 20678;
	#10 counter$count = 20679;
	#10 counter$count = 20680;
	#10 counter$count = 20681;
	#10 counter$count = 20682;
	#10 counter$count = 20683;
	#10 counter$count = 20684;
	#10 counter$count = 20685;
	#10 counter$count = 20686;
	#10 counter$count = 20687;
	#10 counter$count = 20688;
	#10 counter$count = 20689;
	#10 counter$count = 20690;
	#10 counter$count = 20691;
	#10 counter$count = 20692;
	#10 counter$count = 20693;
	#10 counter$count = 20694;
	#10 counter$count = 20695;
	#10 counter$count = 20696;
	#10 counter$count = 20697;
	#10 counter$count = 20698;
	#10 counter$count = 20699;
	#10 counter$count = 20700;
	#10 counter$count = 20701;
	#10 counter$count = 20702;
	#10 counter$count = 20703;
	#10 counter$count = 20704;
	#10 counter$count = 20705;
	#10 counter$count = 20706;
	#10 counter$count = 20707;
	#10 counter$count = 20708;
	#10 counter$count = 20709;
	#10 counter$count = 20710;
	#10 counter$count = 20711;
	#10 counter$count = 20712;
	#10 counter$count = 20713;
	#10 counter$count = 20714;
	#10 counter$count = 20715;
	#10 counter$count = 20716;
	#10 counter$count = 20717;
	#10 counter$count = 20718;
	#10 counter$count = 20719;
	#10 counter$count = 20720;
	#10 counter$count = 20721;
	#10 counter$count = 20722;
	#10 counter$count = 20723;
	#10 counter$count = 20724;
	#10 counter$count = 20725;
	#10 counter$count = 20726;
	#10 counter$count = 20727;
	#10 counter$count = 20728;
	#10 counter$count = 20729;
	#10 counter$count = 20730;
	#10 counter$count = 20731;
	#10 counter$count = 20732;
	#10 counter$count = 20733;
	#10 counter$count = 20734;
	#10 counter$count = 20735;
	#10 counter$count = 20736;
	#10 counter$count = 20737;
	#10 counter$count = 20738;
	#10 counter$count = 20739;
	#10 counter$count = 20740;
	#10 counter$count = 20741;
	#10 counter$count = 20742;
	#10 counter$count = 20743;
	#10 counter$count = 20744;
	#10 counter$count = 20745;
	#10 counter$count = 20746;
	#10 counter$count = 20747;
	#10 counter$count = 20748;
	#10 counter$count = 20749;
	#10 counter$count = 20750;
	#10 counter$count = 20751;
	#10 counter$count = 20752;
	#10 counter$count = 20753;
	#10 counter$count = 20754;
	#10 counter$count = 20755;
	#10 counter$count = 20756;
	#10 counter$count = 20757;
	#10 counter$count = 20758;
	#10 counter$count = 20759;
	#10 counter$count = 20760;
	#10 counter$count = 20761;
	#10 counter$count = 20762;
	#10 counter$count = 20763;
	#10 counter$count = 20764;
	#10 counter$count = 20765;
	#10 counter$count = 20766;
	#10 counter$count = 20767;
	#10 counter$count = 20768;
	#10 counter$count = 20769;
	#10 counter$count = 20770;
	#10 counter$count = 20771;
	#10 counter$count = 20772;
	#10 counter$count = 20773;
	#10 counter$count = 20774;
	#10 counter$count = 20775;
	#10 counter$count = 20776;
	#10 counter$count = 20777;
	#10 counter$count = 20778;
	#10 counter$count = 20779;
	#10 counter$count = 20780;
	#10 counter$count = 20781;
	#10 counter$count = 20782;
	#10 counter$count = 20783;
	#10 counter$count = 20784;
	#10 counter$count = 20785;
	#10 counter$count = 20786;
	#10 counter$count = 20787;
	#10 counter$count = 20788;
	#10 counter$count = 20789;
	#10 counter$count = 20790;
	#10 counter$count = 20791;
	#10 counter$count = 20792;
	#10 counter$count = 20793;
	#10 counter$count = 20794;
	#10 counter$count = 20795;
	#10 counter$count = 20796;
	#10 counter$count = 20797;
	#10 counter$count = 20798;
	#10 counter$count = 20799;
	#10 counter$count = 20800;
	#10 counter$count = 20801;
	#10 counter$count = 20802;
	#10 counter$count = 20803;
	#10 counter$count = 20804;
	#10 counter$count = 20805;
	#10 counter$count = 20806;
	#10 counter$count = 20807;
	#10 counter$count = 20808;
	#10 counter$count = 20809;
	#10 counter$count = 20810;
	#10 counter$count = 20811;
	#10 counter$count = 20812;
	#10 counter$count = 20813;
	#10 counter$count = 20814;
	#10 counter$count = 20815;
	#10 counter$count = 20816;
	#10 counter$count = 20817;
	#10 counter$count = 20818;
	#10 counter$count = 20819;
	#10 counter$count = 20820;
	#10 counter$count = 20821;
	#10 counter$count = 20822;
	#10 counter$count = 20823;
	#10 counter$count = 20824;
	#10 counter$count = 20825;
	#10 counter$count = 20826;
	#10 counter$count = 20827;
	#10 counter$count = 20828;
	#10 counter$count = 20829;
	#10 counter$count = 20830;
	#10 counter$count = 20831;
	#10 counter$count = 20832;
	#10 counter$count = 20833;
	#10 counter$count = 20834;
	#10 counter$count = 20835;
	#10 counter$count = 20836;
	#10 counter$count = 20837;
	#10 counter$count = 20838;
	#10 counter$count = 20839;
	#10 counter$count = 20840;
	#10 counter$count = 20841;
	#10 counter$count = 20842;
	#10 counter$count = 20843;
	#10 counter$count = 20844;
	#10 counter$count = 20845;
	#10 counter$count = 20846;
	#10 counter$count = 20847;
	#10 counter$count = 20848;
	#10 counter$count = 20849;
	#10 counter$count = 20850;
	#10 counter$count = 20851;
	#10 counter$count = 20852;
	#10 counter$count = 20853;
	#10 counter$count = 20854;
	#10 counter$count = 20855;
	#10 counter$count = 20856;
	#10 counter$count = 20857;
	#10 counter$count = 20858;
	#10 counter$count = 20859;
	#10 counter$count = 20860;
	#10 counter$count = 20861;
	#10 counter$count = 20862;
	#10 counter$count = 20863;
	#10 counter$count = 20864;
	#10 counter$count = 20865;
	#10 counter$count = 20866;
	#10 counter$count = 20867;
	#10 counter$count = 20868;
	#10 counter$count = 20869;
	#10 counter$count = 20870;
	#10 counter$count = 20871;
	#10 counter$count = 20872;
	#10 counter$count = 20873;
	#10 counter$count = 20874;
	#10 counter$count = 20875;
	#10 counter$count = 20876;
	#10 counter$count = 20877;
	#10 counter$count = 20878;
	#10 counter$count = 20879;
	#10 counter$count = 20880;
	#10 counter$count = 20881;
	#10 counter$count = 20882;
	#10 counter$count = 20883;
	#10 counter$count = 20884;
	#10 counter$count = 20885;
	#10 counter$count = 20886;
	#10 counter$count = 20887;
	#10 counter$count = 20888;
	#10 counter$count = 20889;
	#10 counter$count = 20890;
	#10 counter$count = 20891;
	#10 counter$count = 20892;
	#10 counter$count = 20893;
	#10 counter$count = 20894;
	#10 counter$count = 20895;
	#10 counter$count = 20896;
	#10 counter$count = 20897;
	#10 counter$count = 20898;
	#10 counter$count = 20899;
	#10 counter$count = 20900;
	#10 counter$count = 20901;
	#10 counter$count = 20902;
	#10 counter$count = 20903;
	#10 counter$count = 20904;
	#10 counter$count = 20905;
	#10 counter$count = 20906;
	#10 counter$count = 20907;
	#10 counter$count = 20908;
	#10 counter$count = 20909;
	#10 counter$count = 20910;
	#10 counter$count = 20911;
	#10 counter$count = 20912;
	#10 counter$count = 20913;
	#10 counter$count = 20914;
	#10 counter$count = 20915;
	#10 counter$count = 20916;
	#10 counter$count = 20917;
	#10 counter$count = 20918;
	#10 counter$count = 20919;
	#10 counter$count = 20920;
	#10 counter$count = 20921;
	#10 counter$count = 20922;
	#10 counter$count = 20923;
	#10 counter$count = 20924;
	#10 counter$count = 20925;
	#10 counter$count = 20926;
	#10 counter$count = 20927;
	#10 counter$count = 20928;
	#10 counter$count = 20929;
	#10 counter$count = 20930;
	#10 counter$count = 20931;
	#10 counter$count = 20932;
	#10 counter$count = 20933;
	#10 counter$count = 20934;
	#10 counter$count = 20935;
	#10 counter$count = 20936;
	#10 counter$count = 20937;
	#10 counter$count = 20938;
	#10 counter$count = 20939;
	#10 counter$count = 20940;
	#10 counter$count = 20941;
	#10 counter$count = 20942;
	#10 counter$count = 20943;
	#10 counter$count = 20944;
	#10 counter$count = 20945;
	#10 counter$count = 20946;
	#10 counter$count = 20947;
	#10 counter$count = 20948;
	#10 counter$count = 20949;
	#10 counter$count = 20950;
	#10 counter$count = 20951;
	#10 counter$count = 20952;
	#10 counter$count = 20953;
	#10 counter$count = 20954;
	#10 counter$count = 20955;
	#10 counter$count = 20956;
	#10 counter$count = 20957;
	#10 counter$count = 20958;
	#10 counter$count = 20959;
	#10 counter$count = 20960;
	#10 counter$count = 20961;
	#10 counter$count = 20962;
	#10 counter$count = 20963;
	#10 counter$count = 20964;
	#10 counter$count = 20965;
	#10 counter$count = 20966;
	#10 counter$count = 20967;
	#10 counter$count = 20968;
	#10 counter$count = 20969;
	#10 counter$count = 20970;
	#10 counter$count = 20971;
	#10 counter$count = 20972;
	#10 counter$count = 20973;
	#10 counter$count = 20974;
	#10 counter$count = 20975;
	#10 counter$count = 20976;
	#10 counter$count = 20977;
	#10 counter$count = 20978;
	#10 counter$count = 20979;
	#10 counter$count = 20980;
	#10 counter$count = 20981;
	#10 counter$count = 20982;
	#10 counter$count = 20983;
	#10 counter$count = 20984;
	#10 counter$count = 20985;
	#10 counter$count = 20986;
	#10 counter$count = 20987;
	#10 counter$count = 20988;
	#10 counter$count = 20989;
	#10 counter$count = 20990;
	#10 counter$count = 20991;
	#10 counter$count = 20992;
	#10 counter$count = 20993;
	#10 counter$count = 20994;
	#10 counter$count = 20995;
	#10 counter$count = 20996;
	#10 counter$count = 20997;
	#10 counter$count = 20998;
	#10 counter$count = 20999;
	#10 counter$count = 21000;
	#10 counter$count = 21001;
	#10 counter$count = 21002;
	#10 counter$count = 21003;
	#10 counter$count = 21004;
	#10 counter$count = 21005;
	#10 counter$count = 21006;
	#10 counter$count = 21007;
	#10 counter$count = 21008;
	#10 counter$count = 21009;
	#10 counter$count = 21010;
	#10 counter$count = 21011;
	#10 counter$count = 21012;
	#10 counter$count = 21013;
	#10 counter$count = 21014;
	#10 counter$count = 21015;
	#10 counter$count = 21016;
	#10 counter$count = 21017;
	#10 counter$count = 21018;
	#10 counter$count = 21019;
	#10 counter$count = 21020;
	#10 counter$count = 21021;
	#10 counter$count = 21022;
	#10 counter$count = 21023;
	#10 counter$count = 21024;
	#10 counter$count = 21025;
	#10 counter$count = 21026;
	#10 counter$count = 21027;
	#10 counter$count = 21028;
	#10 counter$count = 21029;
	#10 counter$count = 21030;
	#10 counter$count = 21031;
	#10 counter$count = 21032;
	#10 counter$count = 21033;
	#10 counter$count = 21034;
	#10 counter$count = 21035;
	#10 counter$count = 21036;
	#10 counter$count = 21037;
	#10 counter$count = 21038;
	#10 counter$count = 21039;
	#10 counter$count = 21040;
	#10 counter$count = 21041;
	#10 counter$count = 21042;
	#10 counter$count = 21043;
	#10 counter$count = 21044;
	#10 counter$count = 21045;
	#10 counter$count = 21046;
	#10 counter$count = 21047;
	#10 counter$count = 21048;
	#10 counter$count = 21049;
	#10 counter$count = 21050;
	#10 counter$count = 21051;
	#10 counter$count = 21052;
	#10 counter$count = 21053;
	#10 counter$count = 21054;
	#10 counter$count = 21055;
	#10 counter$count = 21056;
	#10 counter$count = 21057;
	#10 counter$count = 21058;
	#10 counter$count = 21059;
	#10 counter$count = 21060;
	#10 counter$count = 21061;
	#10 counter$count = 21062;
	#10 counter$count = 21063;
	#10 counter$count = 21064;
	#10 counter$count = 21065;
	#10 counter$count = 21066;
	#10 counter$count = 21067;
	#10 counter$count = 21068;
	#10 counter$count = 21069;
	#10 counter$count = 21070;
	#10 counter$count = 21071;
	#10 counter$count = 21072;
	#10 counter$count = 21073;
	#10 counter$count = 21074;
	#10 counter$count = 21075;
	#10 counter$count = 21076;
	#10 counter$count = 21077;
	#10 counter$count = 21078;
	#10 counter$count = 21079;
	#10 counter$count = 21080;
	#10 counter$count = 21081;
	#10 counter$count = 21082;
	#10 counter$count = 21083;
	#10 counter$count = 21084;
	#10 counter$count = 21085;
	#10 counter$count = 21086;
	#10 counter$count = 21087;
	#10 counter$count = 21088;
	#10 counter$count = 21089;
	#10 counter$count = 21090;
	#10 counter$count = 21091;
	#10 counter$count = 21092;
	#10 counter$count = 21093;
	#10 counter$count = 21094;
	#10 counter$count = 21095;
	#10 counter$count = 21096;
	#10 counter$count = 21097;
	#10 counter$count = 21098;
	#10 counter$count = 21099;
	#10 counter$count = 21100;
	#10 counter$count = 21101;
	#10 counter$count = 21102;
	#10 counter$count = 21103;
	#10 counter$count = 21104;
	#10 counter$count = 21105;
	#10 counter$count = 21106;
	#10 counter$count = 21107;
	#10 counter$count = 21108;
	#10 counter$count = 21109;
	#10 counter$count = 21110;
	#10 counter$count = 21111;
	#10 counter$count = 21112;
	#10 counter$count = 21113;
	#10 counter$count = 21114;
	#10 counter$count = 21115;
	#10 counter$count = 21116;
	#10 counter$count = 21117;
	#10 counter$count = 21118;
	#10 counter$count = 21119;
	#10 counter$count = 21120;
	#10 counter$count = 21121;
	#10 counter$count = 21122;
	#10 counter$count = 21123;
	#10 counter$count = 21124;
	#10 counter$count = 21125;
	#10 counter$count = 21126;
	#10 counter$count = 21127;
	#10 counter$count = 21128;
	#10 counter$count = 21129;
	#10 counter$count = 21130;
	#10 counter$count = 21131;
	#10 counter$count = 21132;
	#10 counter$count = 21133;
	#10 counter$count = 21134;
	#10 counter$count = 21135;
	#10 counter$count = 21136;
	#10 counter$count = 21137;
	#10 counter$count = 21138;
	#10 counter$count = 21139;
	#10 counter$count = 21140;
	#10 counter$count = 21141;
	#10 counter$count = 21142;
	#10 counter$count = 21143;
	#10 counter$count = 21144;
	#10 counter$count = 21145;
	#10 counter$count = 21146;
	#10 counter$count = 21147;
	#10 counter$count = 21148;
	#10 counter$count = 21149;
	#10 counter$count = 21150;
	#10 counter$count = 21151;
	#10 counter$count = 21152;
	#10 counter$count = 21153;
	#10 counter$count = 21154;
	#10 counter$count = 21155;
	#10 counter$count = 21156;
	#10 counter$count = 21157;
	#10 counter$count = 21158;
	#10 counter$count = 21159;
	#10 counter$count = 21160;
	#10 counter$count = 21161;
	#10 counter$count = 21162;
	#10 counter$count = 21163;
	#10 counter$count = 21164;
	#10 counter$count = 21165;
	#10 counter$count = 21166;
	#10 counter$count = 21167;
	#10 counter$count = 21168;
	#10 counter$count = 21169;
	#10 counter$count = 21170;
	#10 counter$count = 21171;
	#10 counter$count = 21172;
	#10 counter$count = 21173;
	#10 counter$count = 21174;
	#10 counter$count = 21175;
	#10 counter$count = 21176;
	#10 counter$count = 21177;
	#10 counter$count = 21178;
	#10 counter$count = 21179;
	#10 counter$count = 21180;
	#10 counter$count = 21181;
	#10 counter$count = 21182;
	#10 counter$count = 21183;
	#10 counter$count = 21184;
	#10 counter$count = 21185;
	#10 counter$count = 21186;
	#10 counter$count = 21187;
	#10 counter$count = 21188;
	#10 counter$count = 21189;
	#10 counter$count = 21190;
	#10 counter$count = 21191;
	#10 counter$count = 21192;
	#10 counter$count = 21193;
	#10 counter$count = 21194;
	#10 counter$count = 21195;
	#10 counter$count = 21196;
	#10 counter$count = 21197;
	#10 counter$count = 21198;
	#10 counter$count = 21199;
	#10 counter$count = 21200;
	#10 counter$count = 21201;
	#10 counter$count = 21202;
	#10 counter$count = 21203;
	#10 counter$count = 21204;
	#10 counter$count = 21205;
	#10 counter$count = 21206;
	#10 counter$count = 21207;
	#10 counter$count = 21208;
	#10 counter$count = 21209;
	#10 counter$count = 21210;
	#10 counter$count = 21211;
	#10 counter$count = 21212;
	#10 counter$count = 21213;
	#10 counter$count = 21214;
	#10 counter$count = 21215;
	#10 counter$count = 21216;
	#10 counter$count = 21217;
	#10 counter$count = 21218;
	#10 counter$count = 21219;
	#10 counter$count = 21220;
	#10 counter$count = 21221;
	#10 counter$count = 21222;
	#10 counter$count = 21223;
	#10 counter$count = 21224;
	#10 counter$count = 21225;
	#10 counter$count = 21226;
	#10 counter$count = 21227;
	#10 counter$count = 21228;
	#10 counter$count = 21229;
	#10 counter$count = 21230;
	#10 counter$count = 21231;
	#10 counter$count = 21232;
	#10 counter$count = 21233;
	#10 counter$count = 21234;
	#10 counter$count = 21235;
	#10 counter$count = 21236;
	#10 counter$count = 21237;
	#10 counter$count = 21238;
	#10 counter$count = 21239;
	#10 counter$count = 21240;
	#10 counter$count = 21241;
	#10 counter$count = 21242;
	#10 counter$count = 21243;
	#10 counter$count = 21244;
	#10 counter$count = 21245;
	#10 counter$count = 21246;
	#10 counter$count = 21247;
	#10 counter$count = 21248;
	#10 counter$count = 21249;
	#10 counter$count = 21250;
	#10 counter$count = 21251;
	#10 counter$count = 21252;
	#10 counter$count = 21253;
	#10 counter$count = 21254;
	#10 counter$count = 21255;
	#10 counter$count = 21256;
	#10 counter$count = 21257;
	#10 counter$count = 21258;
	#10 counter$count = 21259;
	#10 counter$count = 21260;
	#10 counter$count = 21261;
	#10 counter$count = 21262;
	#10 counter$count = 21263;
	#10 counter$count = 21264;
	#10 counter$count = 21265;
	#10 counter$count = 21266;
	#10 counter$count = 21267;
	#10 counter$count = 21268;
	#10 counter$count = 21269;
	#10 counter$count = 21270;
	#10 counter$count = 21271;
	#10 counter$count = 21272;
	#10 counter$count = 21273;
	#10 counter$count = 21274;
	#10 counter$count = 21275;
	#10 counter$count = 21276;
	#10 counter$count = 21277;
	#10 counter$count = 21278;
	#10 counter$count = 21279;
	#10 counter$count = 21280;
	#10 counter$count = 21281;
	#10 counter$count = 21282;
	#10 counter$count = 21283;
	#10 counter$count = 21284;
	#10 counter$count = 21285;
	#10 counter$count = 21286;
	#10 counter$count = 21287;
	#10 counter$count = 21288;
	#10 counter$count = 21289;
	#10 counter$count = 21290;
	#10 counter$count = 21291;
	#10 counter$count = 21292;
	#10 counter$count = 21293;
	#10 counter$count = 21294;
	#10 counter$count = 21295;
	#10 counter$count = 21296;
	#10 counter$count = 21297;
	#10 counter$count = 21298;
	#10 counter$count = 21299;
	#10 counter$count = 21300;
	#10 counter$count = 21301;
	#10 counter$count = 21302;
	#10 counter$count = 21303;
	#10 counter$count = 21304;
	#10 counter$count = 21305;
	#10 counter$count = 21306;
	#10 counter$count = 21307;
	#10 counter$count = 21308;
	#10 counter$count = 21309;
	#10 counter$count = 21310;
	#10 counter$count = 21311;
	#10 counter$count = 21312;
	#10 counter$count = 21313;
	#10 counter$count = 21314;
	#10 counter$count = 21315;
	#10 counter$count = 21316;
	#10 counter$count = 21317;
	#10 counter$count = 21318;
	#10 counter$count = 21319;
	#10 counter$count = 21320;
	#10 counter$count = 21321;
	#10 counter$count = 21322;
	#10 counter$count = 21323;
	#10 counter$count = 21324;
	#10 counter$count = 21325;
	#10 counter$count = 21326;
	#10 counter$count = 21327;
	#10 counter$count = 21328;
	#10 counter$count = 21329;
	#10 counter$count = 21330;
	#10 counter$count = 21331;
	#10 counter$count = 21332;
	#10 counter$count = 21333;
	#10 counter$count = 21334;
	#10 counter$count = 21335;
	#10 counter$count = 21336;
	#10 counter$count = 21337;
	#10 counter$count = 21338;
	#10 counter$count = 21339;
	#10 counter$count = 21340;
	#10 counter$count = 21341;
	#10 counter$count = 21342;
	#10 counter$count = 21343;
	#10 counter$count = 21344;
	#10 counter$count = 21345;
	#10 counter$count = 21346;
	#10 counter$count = 21347;
	#10 counter$count = 21348;
	#10 counter$count = 21349;
	#10 counter$count = 21350;
	#10 counter$count = 21351;
	#10 counter$count = 21352;
	#10 counter$count = 21353;
	#10 counter$count = 21354;
	#10 counter$count = 21355;
	#10 counter$count = 21356;
	#10 counter$count = 21357;
	#10 counter$count = 21358;
	#10 counter$count = 21359;
	#10 counter$count = 21360;
	#10 counter$count = 21361;
	#10 counter$count = 21362;
	#10 counter$count = 21363;
	#10 counter$count = 21364;
	#10 counter$count = 21365;
	#10 counter$count = 21366;
	#10 counter$count = 21367;
	#10 counter$count = 21368;
	#10 counter$count = 21369;
	#10 counter$count = 21370;
	#10 counter$count = 21371;
	#10 counter$count = 21372;
	#10 counter$count = 21373;
	#10 counter$count = 21374;
	#10 counter$count = 21375;
	#10 counter$count = 21376;
	#10 counter$count = 21377;
	#10 counter$count = 21378;
	#10 counter$count = 21379;
	#10 counter$count = 21380;
	#10 counter$count = 21381;
	#10 counter$count = 21382;
	#10 counter$count = 21383;
	#10 counter$count = 21384;
	#10 counter$count = 21385;
	#10 counter$count = 21386;
	#10 counter$count = 21387;
	#10 counter$count = 21388;
	#10 counter$count = 21389;
	#10 counter$count = 21390;
	#10 counter$count = 21391;
	#10 counter$count = 21392;
	#10 counter$count = 21393;
	#10 counter$count = 21394;
	#10 counter$count = 21395;
	#10 counter$count = 21396;
	#10 counter$count = 21397;
	#10 counter$count = 21398;
	#10 counter$count = 21399;
	#10 counter$count = 21400;
	#10 counter$count = 21401;
	#10 counter$count = 21402;
	#10 counter$count = 21403;
	#10 counter$count = 21404;
	#10 counter$count = 21405;
	#10 counter$count = 21406;
	#10 counter$count = 21407;
	#10 counter$count = 21408;
	#10 counter$count = 21409;
	#10 counter$count = 21410;
	#10 counter$count = 21411;
	#10 counter$count = 21412;
	#10 counter$count = 21413;
	#10 counter$count = 21414;
	#10 counter$count = 21415;
	#10 counter$count = 21416;
	#10 counter$count = 21417;
	#10 counter$count = 21418;
	#10 counter$count = 21419;
	#10 counter$count = 21420;
	#10 counter$count = 21421;
	#10 counter$count = 21422;
	#10 counter$count = 21423;
	#10 counter$count = 21424;
	#10 counter$count = 21425;
	#10 counter$count = 21426;
	#10 counter$count = 21427;
	#10 counter$count = 21428;
	#10 counter$count = 21429;
	#10 counter$count = 21430;
	#10 counter$count = 21431;
	#10 counter$count = 21432;
	#10 counter$count = 21433;
	#10 counter$count = 21434;
	#10 counter$count = 21435;
	#10 counter$count = 21436;
	#10 counter$count = 21437;
	#10 counter$count = 21438;
	#10 counter$count = 21439;
	#10 counter$count = 21440;
	#10 counter$count = 21441;
	#10 counter$count = 21442;
	#10 counter$count = 21443;
	#10 counter$count = 21444;
	#10 counter$count = 21445;
	#10 counter$count = 21446;
	#10 counter$count = 21447;
	#10 counter$count = 21448;
	#10 counter$count = 21449;
	#10 counter$count = 21450;
	#10 counter$count = 21451;
	#10 counter$count = 21452;
	#10 counter$count = 21453;
	#10 counter$count = 21454;
	#10 counter$count = 21455;
	#10 counter$count = 21456;
	#10 counter$count = 21457;
	#10 counter$count = 21458;
	#10 counter$count = 21459;
	#10 counter$count = 21460;
	#10 counter$count = 21461;
	#10 counter$count = 21462;
	#10 counter$count = 21463;
	#10 counter$count = 21464;
	#10 counter$count = 21465;
	#10 counter$count = 21466;
	#10 counter$count = 21467;
	#10 counter$count = 21468;
	#10 counter$count = 21469;
	#10 counter$count = 21470;
	#10 counter$count = 21471;
	#10 counter$count = 21472;
	#10 counter$count = 21473;
	#10 counter$count = 21474;
	#10 counter$count = 21475;
	#10 counter$count = 21476;
	#10 counter$count = 21477;
	#10 counter$count = 21478;
	#10 counter$count = 21479;
	#10 counter$count = 21480;
	#10 counter$count = 21481;
	#10 counter$count = 21482;
	#10 counter$count = 21483;
	#10 counter$count = 21484;
	#10 counter$count = 21485;
	#10 counter$count = 21486;
	#10 counter$count = 21487;
	#10 counter$count = 21488;
	#10 counter$count = 21489;
	#10 counter$count = 21490;
	#10 counter$count = 21491;
	#10 counter$count = 21492;
	#10 counter$count = 21493;
	#10 counter$count = 21494;
	#10 counter$count = 21495;
	#10 counter$count = 21496;
	#10 counter$count = 21497;
	#10 counter$count = 21498;
	#10 counter$count = 21499;
	#10 counter$count = 21500;
	#10 counter$count = 21501;
	#10 counter$count = 21502;
	#10 counter$count = 21503;
	#10 counter$count = 21504;
	#10 counter$count = 21505;
	#10 counter$count = 21506;
	#10 counter$count = 21507;
	#10 counter$count = 21508;
	#10 counter$count = 21509;
	#10 counter$count = 21510;
	#10 counter$count = 21511;
	#10 counter$count = 21512;
	#10 counter$count = 21513;
	#10 counter$count = 21514;
	#10 counter$count = 21515;
	#10 counter$count = 21516;
	#10 counter$count = 21517;
	#10 counter$count = 21518;
	#10 counter$count = 21519;
	#10 counter$count = 21520;
	#10 counter$count = 21521;
	#10 counter$count = 21522;
	#10 counter$count = 21523;
	#10 counter$count = 21524;
	#10 counter$count = 21525;
	#10 counter$count = 21526;
	#10 counter$count = 21527;
	#10 counter$count = 21528;
	#10 counter$count = 21529;
	#10 counter$count = 21530;
	#10 counter$count = 21531;
	#10 counter$count = 21532;
	#10 counter$count = 21533;
	#10 counter$count = 21534;
	#10 counter$count = 21535;
	#10 counter$count = 21536;
	#10 counter$count = 21537;
	#10 counter$count = 21538;
	#10 counter$count = 21539;
	#10 counter$count = 21540;
	#10 counter$count = 21541;
	#10 counter$count = 21542;
	#10 counter$count = 21543;
	#10 counter$count = 21544;
	#10 counter$count = 21545;
	#10 counter$count = 21546;
	#10 counter$count = 21547;
	#10 counter$count = 21548;
	#10 counter$count = 21549;
	#10 counter$count = 21550;
	#10 counter$count = 21551;
	#10 counter$count = 21552;
	#10 counter$count = 21553;
	#10 counter$count = 21554;
	#10 counter$count = 21555;
	#10 counter$count = 21556;
	#10 counter$count = 21557;
	#10 counter$count = 21558;
	#10 counter$count = 21559;
	#10 counter$count = 21560;
	#10 counter$count = 21561;
	#10 counter$count = 21562;
	#10 counter$count = 21563;
	#10 counter$count = 21564;
	#10 counter$count = 21565;
	#10 counter$count = 21566;
	#10 counter$count = 21567;
	#10 counter$count = 21568;
	#10 counter$count = 21569;
	#10 counter$count = 21570;
	#10 counter$count = 21571;
	#10 counter$count = 21572;
	#10 counter$count = 21573;
	#10 counter$count = 21574;
	#10 counter$count = 21575;
	#10 counter$count = 21576;
	#10 counter$count = 21577;
	#10 counter$count = 21578;
	#10 counter$count = 21579;
	#10 counter$count = 21580;
	#10 counter$count = 21581;
	#10 counter$count = 21582;
	#10 counter$count = 21583;
	#10 counter$count = 21584;
	#10 counter$count = 21585;
	#10 counter$count = 21586;
	#10 counter$count = 21587;
	#10 counter$count = 21588;
	#10 counter$count = 21589;
	#10 counter$count = 21590;
	#10 counter$count = 21591;
	#10 counter$count = 21592;
	#10 counter$count = 21593;
	#10 counter$count = 21594;
	#10 counter$count = 21595;
	#10 counter$count = 21596;
	#10 counter$count = 21597;
	#10 counter$count = 21598;
	#10 counter$count = 21599;
	#10 counter$count = 21600;
	#10 counter$count = 21601;
	#10 counter$count = 21602;
	#10 counter$count = 21603;
	#10 counter$count = 21604;
	#10 counter$count = 21605;
	#10 counter$count = 21606;
	#10 counter$count = 21607;
	#10 counter$count = 21608;
	#10 counter$count = 21609;
	#10 counter$count = 21610;
	#10 counter$count = 21611;
	#10 counter$count = 21612;
	#10 counter$count = 21613;
	#10 counter$count = 21614;
	#10 counter$count = 21615;
	#10 counter$count = 21616;
	#10 counter$count = 21617;
	#10 counter$count = 21618;
	#10 counter$count = 21619;
	#10 counter$count = 21620;
	#10 counter$count = 21621;
	#10 counter$count = 21622;
	#10 counter$count = 21623;
	#10 counter$count = 21624;
	#10 counter$count = 21625;
	#10 counter$count = 21626;
	#10 counter$count = 21627;
	#10 counter$count = 21628;
	#10 counter$count = 21629;
	#10 counter$count = 21630;
	#10 counter$count = 21631;
	#10 counter$count = 21632;
	#10 counter$count = 21633;
	#10 counter$count = 21634;
	#10 counter$count = 21635;
	#10 counter$count = 21636;
	#10 counter$count = 21637;
	#10 counter$count = 21638;
	#10 counter$count = 21639;
	#10 counter$count = 21640;
	#10 counter$count = 21641;
	#10 counter$count = 21642;
	#10 counter$count = 21643;
	#10 counter$count = 21644;
	#10 counter$count = 21645;
	#10 counter$count = 21646;
	#10 counter$count = 21647;
	#10 counter$count = 21648;
	#10 counter$count = 21649;
	#10 counter$count = 21650;
	#10 counter$count = 21651;
	#10 counter$count = 21652;
	#10 counter$count = 21653;
	#10 counter$count = 21654;
	#10 counter$count = 21655;
	#10 counter$count = 21656;
	#10 counter$count = 21657;
	#10 counter$count = 21658;
	#10 counter$count = 21659;
	#10 counter$count = 21660;
	#10 counter$count = 21661;
	#10 counter$count = 21662;
	#10 counter$count = 21663;
	#10 counter$count = 21664;
	#10 counter$count = 21665;
	#10 counter$count = 21666;
	#10 counter$count = 21667;
	#10 counter$count = 21668;
	#10 counter$count = 21669;
	#10 counter$count = 21670;
	#10 counter$count = 21671;
	#10 counter$count = 21672;
	#10 counter$count = 21673;
	#10 counter$count = 21674;
	#10 counter$count = 21675;
	#10 counter$count = 21676;
	#10 counter$count = 21677;
	#10 counter$count = 21678;
	#10 counter$count = 21679;
	#10 counter$count = 21680;
	#10 counter$count = 21681;
	#10 counter$count = 21682;
	#10 counter$count = 21683;
	#10 counter$count = 21684;
	#10 counter$count = 21685;
	#10 counter$count = 21686;
	#10 counter$count = 21687;
	#10 counter$count = 21688;
	#10 counter$count = 21689;
	#10 counter$count = 21690;
	#10 counter$count = 21691;
	#10 counter$count = 21692;
	#10 counter$count = 21693;
	#10 counter$count = 21694;
	#10 counter$count = 21695;
	#10 counter$count = 21696;
	#10 counter$count = 21697;
	#10 counter$count = 21698;
	#10 counter$count = 21699;
	#10 counter$count = 21700;
	#10 counter$count = 21701;
	#10 counter$count = 21702;
	#10 counter$count = 21703;
	#10 counter$count = 21704;
	#10 counter$count = 21705;
	#10 counter$count = 21706;
	#10 counter$count = 21707;
	#10 counter$count = 21708;
	#10 counter$count = 21709;
	#10 counter$count = 21710;
	#10 counter$count = 21711;
	#10 counter$count = 21712;
	#10 counter$count = 21713;
	#10 counter$count = 21714;
	#10 counter$count = 21715;
	#10 counter$count = 21716;
	#10 counter$count = 21717;
	#10 counter$count = 21718;
	#10 counter$count = 21719;
	#10 counter$count = 21720;
	#10 counter$count = 21721;
	#10 counter$count = 21722;
	#10 counter$count = 21723;
	#10 counter$count = 21724;
	#10 counter$count = 21725;
	#10 counter$count = 21726;
	#10 counter$count = 21727;
	#10 counter$count = 21728;
	#10 counter$count = 21729;
	#10 counter$count = 21730;
	#10 counter$count = 21731;
	#10 counter$count = 21732;
	#10 counter$count = 21733;
	#10 counter$count = 21734;
	#10 counter$count = 21735;
	#10 counter$count = 21736;
	#10 counter$count = 21737;
	#10 counter$count = 21738;
	#10 counter$count = 21739;
	#10 counter$count = 21740;
	#10 counter$count = 21741;
	#10 counter$count = 21742;
	#10 counter$count = 21743;
	#10 counter$count = 21744;
	#10 counter$count = 21745;
	#10 counter$count = 21746;
	#10 counter$count = 21747;
	#10 counter$count = 21748;
	#10 counter$count = 21749;
	#10 counter$count = 21750;
	#10 counter$count = 21751;
	#10 counter$count = 21752;
	#10 counter$count = 21753;
	#10 counter$count = 21754;
	#10 counter$count = 21755;
	#10 counter$count = 21756;
	#10 counter$count = 21757;
	#10 counter$count = 21758;
	#10 counter$count = 21759;
	#10 counter$count = 21760;
	#10 counter$count = 21761;
	#10 counter$count = 21762;
	#10 counter$count = 21763;
	#10 counter$count = 21764;
	#10 counter$count = 21765;
	#10 counter$count = 21766;
	#10 counter$count = 21767;
	#10 counter$count = 21768;
	#10 counter$count = 21769;
	#10 counter$count = 21770;
	#10 counter$count = 21771;
	#10 counter$count = 21772;
	#10 counter$count = 21773;
	#10 counter$count = 21774;
	#10 counter$count = 21775;
	#10 counter$count = 21776;
	#10 counter$count = 21777;
	#10 counter$count = 21778;
	#10 counter$count = 21779;
	#10 counter$count = 21780;
	#10 counter$count = 21781;
	#10 counter$count = 21782;
	#10 counter$count = 21783;
	#10 counter$count = 21784;
	#10 counter$count = 21785;
	#10 counter$count = 21786;
	#10 counter$count = 21787;
	#10 counter$count = 21788;
	#10 counter$count = 21789;
	#10 counter$count = 21790;
	#10 counter$count = 21791;
	#10 counter$count = 21792;
	#10 counter$count = 21793;
	#10 counter$count = 21794;
	#10 counter$count = 21795;
	#10 counter$count = 21796;
	#10 counter$count = 21797;
	#10 counter$count = 21798;
	#10 counter$count = 21799;
	#10 counter$count = 21800;
	#10 counter$count = 21801;
	#10 counter$count = 21802;
	#10 counter$count = 21803;
	#10 counter$count = 21804;
	#10 counter$count = 21805;
	#10 counter$count = 21806;
	#10 counter$count = 21807;
	#10 counter$count = 21808;
	#10 counter$count = 21809;
	#10 counter$count = 21810;
	#10 counter$count = 21811;
	#10 counter$count = 21812;
	#10 counter$count = 21813;
	#10 counter$count = 21814;
	#10 counter$count = 21815;
	#10 counter$count = 21816;
	#10 counter$count = 21817;
	#10 counter$count = 21818;
	#10 counter$count = 21819;
	#10 counter$count = 21820;
	#10 counter$count = 21821;
	#10 counter$count = 21822;
	#10 counter$count = 21823;
	#10 counter$count = 21824;
	#10 counter$count = 21825;
	#10 counter$count = 21826;
	#10 counter$count = 21827;
	#10 counter$count = 21828;
	#10 counter$count = 21829;
	#10 counter$count = 21830;
	#10 counter$count = 21831;
	#10 counter$count = 21832;
	#10 counter$count = 21833;
	#10 counter$count = 21834;
	#10 counter$count = 21835;
	#10 counter$count = 21836;
	#10 counter$count = 21837;
	#10 counter$count = 21838;
	#10 counter$count = 21839;
	#10 counter$count = 21840;
	#10 counter$count = 21841;
	#10 counter$count = 21842;
	#10 counter$count = 21843;
	#10 counter$count = 21844;
	#10 counter$count = 21845;
	#10 counter$count = 21846;
	#10 counter$count = 21847;
	#10 counter$count = 21848;
	#10 counter$count = 21849;
	#10 counter$count = 21850;
	#10 counter$count = 21851;
	#10 counter$count = 21852;
	#10 counter$count = 21853;
	#10 counter$count = 21854;
	#10 counter$count = 21855;
	#10 counter$count = 21856;
	#10 counter$count = 21857;
	#10 counter$count = 21858;
	#10 counter$count = 21859;
	#10 counter$count = 21860;
	#10 counter$count = 21861;
	#10 counter$count = 21862;
	#10 counter$count = 21863;
	#10 counter$count = 21864;
	#10 counter$count = 21865;
	#10 counter$count = 21866;
	#10 counter$count = 21867;
	#10 counter$count = 21868;
	#10 counter$count = 21869;
	#10 counter$count = 21870;
	#10 counter$count = 21871;
	#10 counter$count = 21872;
	#10 counter$count = 21873;
	#10 counter$count = 21874;
	#10 counter$count = 21875;
	#10 counter$count = 21876;
	#10 counter$count = 21877;
	#10 counter$count = 21878;
	#10 counter$count = 21879;
	#10 counter$count = 21880;
	#10 counter$count = 21881;
	#10 counter$count = 21882;
	#10 counter$count = 21883;
	#10 counter$count = 21884;
	#10 counter$count = 21885;
	#10 counter$count = 21886;
	#10 counter$count = 21887;
	#10 counter$count = 21888;
	#10 counter$count = 21889;
	#10 counter$count = 21890;
	#10 counter$count = 21891;
	#10 counter$count = 21892;
	#10 counter$count = 21893;
	#10 counter$count = 21894;
	#10 counter$count = 21895;
	#10 counter$count = 21896;
	#10 counter$count = 21897;
	#10 counter$count = 21898;
	#10 counter$count = 21899;
	#10 counter$count = 21900;
	#10 counter$count = 21901;
	#10 counter$count = 21902;
	#10 counter$count = 21903;
	#10 counter$count = 21904;
	#10 counter$count = 21905;
	#10 counter$count = 21906;
	#10 counter$count = 21907;
	#10 counter$count = 21908;
	#10 counter$count = 21909;
	#10 counter$count = 21910;
	#10 counter$count = 21911;
	#10 counter$count = 21912;
	#10 counter$count = 21913;
	#10 counter$count = 21914;
	#10 counter$count = 21915;
	#10 counter$count = 21916;
	#10 counter$count = 21917;
	#10 counter$count = 21918;
	#10 counter$count = 21919;
	#10 counter$count = 21920;
	#10 counter$count = 21921;
	#10 counter$count = 21922;
	#10 counter$count = 21923;
	#10 counter$count = 21924;
	#10 counter$count = 21925;
	#10 counter$count = 21926;
	#10 counter$count = 21927;
	#10 counter$count = 21928;
	#10 counter$count = 21929;
	#10 counter$count = 21930;
	#10 counter$count = 21931;
	#10 counter$count = 21932;
	#10 counter$count = 21933;
	#10 counter$count = 21934;
	#10 counter$count = 21935;
	#10 counter$count = 21936;
	#10 counter$count = 21937;
	#10 counter$count = 21938;
	#10 counter$count = 21939;
	#10 counter$count = 21940;
	#10 counter$count = 21941;
	#10 counter$count = 21942;
	#10 counter$count = 21943;
	#10 counter$count = 21944;
	#10 counter$count = 21945;
	#10 counter$count = 21946;
	#10 counter$count = 21947;
	#10 counter$count = 21948;
	#10 counter$count = 21949;
	#10 counter$count = 21950;
	#10 counter$count = 21951;
	#10 counter$count = 21952;
	#10 counter$count = 21953;
	#10 counter$count = 21954;
	#10 counter$count = 21955;
	#10 counter$count = 21956;
	#10 counter$count = 21957;
	#10 counter$count = 21958;
	#10 counter$count = 21959;
	#10 counter$count = 21960;
	#10 counter$count = 21961;
	#10 counter$count = 21962;
	#10 counter$count = 21963;
	#10 counter$count = 21964;
	#10 counter$count = 21965;
	#10 counter$count = 21966;
	#10 counter$count = 21967;
	#10 counter$count = 21968;
	#10 counter$count = 21969;
	#10 counter$count = 21970;
	#10 counter$count = 21971;
	#10 counter$count = 21972;
	#10 counter$count = 21973;
	#10 counter$count = 21974;
	#10 counter$count = 21975;
	#10 counter$count = 21976;
	#10 counter$count = 21977;
	#10 counter$count = 21978;
	#10 counter$count = 21979;
	#10 counter$count = 21980;
	#10 counter$count = 21981;
	#10 counter$count = 21982;
	#10 counter$count = 21983;
	#10 counter$count = 21984;
	#10 counter$count = 21985;
	#10 counter$count = 21986;
	#10 counter$count = 21987;
	#10 counter$count = 21988;
	#10 counter$count = 21989;
	#10 counter$count = 21990;
	#10 counter$count = 21991;
	#10 counter$count = 21992;
	#10 counter$count = 21993;
	#10 counter$count = 21994;
	#10 counter$count = 21995;
	#10 counter$count = 21996;
	#10 counter$count = 21997;
	#10 counter$count = 21998;
	#10 counter$count = 21999;
	#10 counter$count = 22000;
	#10 counter$count = 22001;
	#10 counter$count = 22002;
	#10 counter$count = 22003;
	#10 counter$count = 22004;
	#10 counter$count = 22005;
	#10 counter$count = 22006;
	#10 counter$count = 22007;
	#10 counter$count = 22008;
	#10 counter$count = 22009;
	#10 counter$count = 22010;
	#10 counter$count = 22011;
	#10 counter$count = 22012;
	#10 counter$count = 22013;
	#10 counter$count = 22014;
	#10 counter$count = 22015;
	#10 counter$count = 22016;
	#10 counter$count = 22017;
	#10 counter$count = 22018;
	#10 counter$count = 22019;
	#10 counter$count = 22020;
	#10 counter$count = 22021;
	#10 counter$count = 22022;
	#10 counter$count = 22023;
	#10 counter$count = 22024;
	#10 counter$count = 22025;
	#10 counter$count = 22026;
	#10 counter$count = 22027;
	#10 counter$count = 22028;
	#10 counter$count = 22029;
	#10 counter$count = 22030;
	#10 counter$count = 22031;
	#10 counter$count = 22032;
	#10 counter$count = 22033;
	#10 counter$count = 22034;
	#10 counter$count = 22035;
	#10 counter$count = 22036;
	#10 counter$count = 22037;
	#10 counter$count = 22038;
	#10 counter$count = 22039;
	#10 counter$count = 22040;
	#10 counter$count = 22041;
	#10 counter$count = 22042;
	#10 counter$count = 22043;
	#10 counter$count = 22044;
	#10 counter$count = 22045;
	#10 counter$count = 22046;
	#10 counter$count = 22047;
	#10 counter$count = 22048;
	#10 counter$count = 22049;
	#10 counter$count = 22050;
	#10 counter$count = 22051;
	#10 counter$count = 22052;
	#10 counter$count = 22053;
	#10 counter$count = 22054;
	#10 counter$count = 22055;
	#10 counter$count = 22056;
	#10 counter$count = 22057;
	#10 counter$count = 22058;
	#10 counter$count = 22059;
	#10 counter$count = 22060;
	#10 counter$count = 22061;
	#10 counter$count = 22062;
	#10 counter$count = 22063;
	#10 counter$count = 22064;
	#10 counter$count = 22065;
	#10 counter$count = 22066;
	#10 counter$count = 22067;
	#10 counter$count = 22068;
	#10 counter$count = 22069;
	#10 counter$count = 22070;
	#10 counter$count = 22071;
	#10 counter$count = 22072;
	#10 counter$count = 22073;
	#10 counter$count = 22074;
	#10 counter$count = 22075;
	#10 counter$count = 22076;
	#10 counter$count = 22077;
	#10 counter$count = 22078;
	#10 counter$count = 22079;
	#10 counter$count = 22080;
	#10 counter$count = 22081;
	#10 counter$count = 22082;
	#10 counter$count = 22083;
	#10 counter$count = 22084;
	#10 counter$count = 22085;
	#10 counter$count = 22086;
	#10 counter$count = 22087;
	#10 counter$count = 22088;
	#10 counter$count = 22089;
	#10 counter$count = 22090;
	#10 counter$count = 22091;
	#10 counter$count = 22092;
	#10 counter$count = 22093;
	#10 counter$count = 22094;
	#10 counter$count = 22095;
	#10 counter$count = 22096;
	#10 counter$count = 22097;
	#10 counter$count = 22098;
	#10 counter$count = 22099;
	#10 counter$count = 22100;
	#10 counter$count = 22101;
	#10 counter$count = 22102;
	#10 counter$count = 22103;
	#10 counter$count = 22104;
	#10 counter$count = 22105;
	#10 counter$count = 22106;
	#10 counter$count = 22107;
	#10 counter$count = 22108;
	#10 counter$count = 22109;
	#10 counter$count = 22110;
	#10 counter$count = 22111;
	#10 counter$count = 22112;
	#10 counter$count = 22113;
	#10 counter$count = 22114;
	#10 counter$count = 22115;
	#10 counter$count = 22116;
	#10 counter$count = 22117;
	#10 counter$count = 22118;
	#10 counter$count = 22119;
	#10 counter$count = 22120;
	#10 counter$count = 22121;
	#10 counter$count = 22122;
	#10 counter$count = 22123;
	#10 counter$count = 22124;
	#10 counter$count = 22125;
	#10 counter$count = 22126;
	#10 counter$count = 22127;
	#10 counter$count = 22128;
	#10 counter$count = 22129;
	#10 counter$count = 22130;
	#10 counter$count = 22131;
	#10 counter$count = 22132;
	#10 counter$count = 22133;
	#10 counter$count = 22134;
	#10 counter$count = 22135;
	#10 counter$count = 22136;
	#10 counter$count = 22137;
	#10 counter$count = 22138;
	#10 counter$count = 22139;
	#10 counter$count = 22140;
	#10 counter$count = 22141;
	#10 counter$count = 22142;
	#10 counter$count = 22143;
	#10 counter$count = 22144;
	#10 counter$count = 22145;
	#10 counter$count = 22146;
	#10 counter$count = 22147;
	#10 counter$count = 22148;
	#10 counter$count = 22149;
	#10 counter$count = 22150;
	#10 counter$count = 22151;
	#10 counter$count = 22152;
	#10 counter$count = 22153;
	#10 counter$count = 22154;
	#10 counter$count = 22155;
	#10 counter$count = 22156;
	#10 counter$count = 22157;
	#10 counter$count = 22158;
	#10 counter$count = 22159;
	#10 counter$count = 22160;
	#10 counter$count = 22161;
	#10 counter$count = 22162;
	#10 counter$count = 22163;
	#10 counter$count = 22164;
	#10 counter$count = 22165;
	#10 counter$count = 22166;
	#10 counter$count = 22167;
	#10 counter$count = 22168;
	#10 counter$count = 22169;
	#10 counter$count = 22170;
	#10 counter$count = 22171;
	#10 counter$count = 22172;
	#10 counter$count = 22173;
	#10 counter$count = 22174;
	#10 counter$count = 22175;
	#10 counter$count = 22176;
	#10 counter$count = 22177;
	#10 counter$count = 22178;
	#10 counter$count = 22179;
	#10 counter$count = 22180;
	#10 counter$count = 22181;
	#10 counter$count = 22182;
	#10 counter$count = 22183;
	#10 counter$count = 22184;
	#10 counter$count = 22185;
	#10 counter$count = 22186;
	#10 counter$count = 22187;
	#10 counter$count = 22188;
	#10 counter$count = 22189;
	#10 counter$count = 22190;
	#10 counter$count = 22191;
	#10 counter$count = 22192;
	#10 counter$count = 22193;
	#10 counter$count = 22194;
	#10 counter$count = 22195;
	#10 counter$count = 22196;
	#10 counter$count = 22197;
	#10 counter$count = 22198;
	#10 counter$count = 22199;
	#10 counter$count = 22200;
	#10 counter$count = 22201;
	#10 counter$count = 22202;
	#10 counter$count = 22203;
	#10 counter$count = 22204;
	#10 counter$count = 22205;
	#10 counter$count = 22206;
	#10 counter$count = 22207;
	#10 counter$count = 22208;
	#10 counter$count = 22209;
	#10 counter$count = 22210;
	#10 counter$count = 22211;
	#10 counter$count = 22212;
	#10 counter$count = 22213;
	#10 counter$count = 22214;
	#10 counter$count = 22215;
	#10 counter$count = 22216;
	#10 counter$count = 22217;
	#10 counter$count = 22218;
	#10 counter$count = 22219;
	#10 counter$count = 22220;
	#10 counter$count = 22221;
	#10 counter$count = 22222;
	#10 counter$count = 22223;
	#10 counter$count = 22224;
	#10 counter$count = 22225;
	#10 counter$count = 22226;
	#10 counter$count = 22227;
	#10 counter$count = 22228;
	#10 counter$count = 22229;
	#10 counter$count = 22230;
	#10 counter$count = 22231;
	#10 counter$count = 22232;
	#10 counter$count = 22233;
	#10 counter$count = 22234;
	#10 counter$count = 22235;
	#10 counter$count = 22236;
	#10 counter$count = 22237;
	#10 counter$count = 22238;
	#10 counter$count = 22239;
	#10 counter$count = 22240;
	#10 counter$count = 22241;
	#10 counter$count = 22242;
	#10 counter$count = 22243;
	#10 counter$count = 22244;
	#10 counter$count = 22245;
	#10 counter$count = 22246;
	#10 counter$count = 22247;
	#10 counter$count = 22248;
	#10 counter$count = 22249;
	#10 counter$count = 22250;
	#10 counter$count = 22251;
	#10 counter$count = 22252;
	#10 counter$count = 22253;
	#10 counter$count = 22254;
	#10 counter$count = 22255;
	#10 counter$count = 22256;
	#10 counter$count = 22257;
	#10 counter$count = 22258;
	#10 counter$count = 22259;
	#10 counter$count = 22260;
	#10 counter$count = 22261;
	#10 counter$count = 22262;
	#10 counter$count = 22263;
	#10 counter$count = 22264;
	#10 counter$count = 22265;
	#10 counter$count = 22266;
	#10 counter$count = 22267;
	#10 counter$count = 22268;
	#10 counter$count = 22269;
	#10 counter$count = 22270;
	#10 counter$count = 22271;
	#10 counter$count = 22272;
	#10 counter$count = 22273;
	#10 counter$count = 22274;
	#10 counter$count = 22275;
	#10 counter$count = 22276;
	#10 counter$count = 22277;
	#10 counter$count = 22278;
	#10 counter$count = 22279;
	#10 counter$count = 22280;
	#10 counter$count = 22281;
	#10 counter$count = 22282;
	#10 counter$count = 22283;
	#10 counter$count = 22284;
	#10 counter$count = 22285;
	#10 counter$count = 22286;
	#10 counter$count = 22287;
	#10 counter$count = 22288;
	#10 counter$count = 22289;
	#10 counter$count = 22290;
	#10 counter$count = 22291;
	#10 counter$count = 22292;
	#10 counter$count = 22293;
	#10 counter$count = 22294;
	#10 counter$count = 22295;
	#10 counter$count = 22296;
	#10 counter$count = 22297;
	#10 counter$count = 22298;
	#10 counter$count = 22299;
	#10 counter$count = 22300;
	#10 counter$count = 22301;
	#10 counter$count = 22302;
	#10 counter$count = 22303;
	#10 counter$count = 22304;
	#10 counter$count = 22305;
	#10 counter$count = 22306;
	#10 counter$count = 22307;
	#10 counter$count = 22308;
	#10 counter$count = 22309;
	#10 counter$count = 22310;
	#10 counter$count = 22311;
	#10 counter$count = 22312;
	#10 counter$count = 22313;
	#10 counter$count = 22314;
	#10 counter$count = 22315;
	#10 counter$count = 22316;
	#10 counter$count = 22317;
	#10 counter$count = 22318;
	#10 counter$count = 22319;
	#10 counter$count = 22320;
	#10 counter$count = 22321;
	#10 counter$count = 22322;
	#10 counter$count = 22323;
	#10 counter$count = 22324;
	#10 counter$count = 22325;
	#10 counter$count = 22326;
	#10 counter$count = 22327;
	#10 counter$count = 22328;
	#10 counter$count = 22329;
	#10 counter$count = 22330;
	#10 counter$count = 22331;
	#10 counter$count = 22332;
	#10 counter$count = 22333;
	#10 counter$count = 22334;
	#10 counter$count = 22335;
	#10 counter$count = 22336;
	#10 counter$count = 22337;
	#10 counter$count = 22338;
	#10 counter$count = 22339;
	#10 counter$count = 22340;
	#10 counter$count = 22341;
	#10 counter$count = 22342;
	#10 counter$count = 22343;
	#10 counter$count = 22344;
	#10 counter$count = 22345;
	#10 counter$count = 22346;
	#10 counter$count = 22347;
	#10 counter$count = 22348;
	#10 counter$count = 22349;
	#10 counter$count = 22350;
	#10 counter$count = 22351;
	#10 counter$count = 22352;
	#10 counter$count = 22353;
	#10 counter$count = 22354;
	#10 counter$count = 22355;
	#10 counter$count = 22356;
	#10 counter$count = 22357;
	#10 counter$count = 22358;
	#10 counter$count = 22359;
	#10 counter$count = 22360;
	#10 counter$count = 22361;
	#10 counter$count = 22362;
	#10 counter$count = 22363;
	#10 counter$count = 22364;
	#10 counter$count = 22365;
	#10 counter$count = 22366;
	#10 counter$count = 22367;
	#10 counter$count = 22368;
	#10 counter$count = 22369;
	#10 counter$count = 22370;
	#10 counter$count = 22371;
	#10 counter$count = 22372;
	#10 counter$count = 22373;
	#10 counter$count = 22374;
	#10 counter$count = 22375;
	#10 counter$count = 22376;
	#10 counter$count = 22377;
	#10 counter$count = 22378;
	#10 counter$count = 22379;
	#10 counter$count = 22380;
	#10 counter$count = 22381;
	#10 counter$count = 22382;
	#10 counter$count = 22383;
	#10 counter$count = 22384;
	#10 counter$count = 22385;
	#10 counter$count = 22386;
	#10 counter$count = 22387;
	#10 counter$count = 22388;
	#10 counter$count = 22389;
	#10 counter$count = 22390;
	#10 counter$count = 22391;
	#10 counter$count = 22392;
	#10 counter$count = 22393;
	#10 counter$count = 22394;
	#10 counter$count = 22395;
	#10 counter$count = 22396;
	#10 counter$count = 22397;
	#10 counter$count = 22398;
	#10 counter$count = 22399;
	#10 counter$count = 22400;
	#10 counter$count = 22401;
	#10 counter$count = 22402;
	#10 counter$count = 22403;
	#10 counter$count = 22404;
	#10 counter$count = 22405;
	#10 counter$count = 22406;
	#10 counter$count = 22407;
	#10 counter$count = 22408;
	#10 counter$count = 22409;
	#10 counter$count = 22410;
	#10 counter$count = 22411;
	#10 counter$count = 22412;
	#10 counter$count = 22413;
	#10 counter$count = 22414;
	#10 counter$count = 22415;
	#10 counter$count = 22416;
	#10 counter$count = 22417;
	#10 counter$count = 22418;
	#10 counter$count = 22419;
	#10 counter$count = 22420;
	#10 counter$count = 22421;
	#10 counter$count = 22422;
	#10 counter$count = 22423;
	#10 counter$count = 22424;
	#10 counter$count = 22425;
	#10 counter$count = 22426;
	#10 counter$count = 22427;
	#10 counter$count = 22428;
	#10 counter$count = 22429;
	#10 counter$count = 22430;
	#10 counter$count = 22431;
	#10 counter$count = 22432;
	#10 counter$count = 22433;
	#10 counter$count = 22434;
	#10 counter$count = 22435;
	#10 counter$count = 22436;
	#10 counter$count = 22437;
	#10 counter$count = 22438;
	#10 counter$count = 22439;
	#10 counter$count = 22440;
	#10 counter$count = 22441;
	#10 counter$count = 22442;
	#10 counter$count = 22443;
	#10 counter$count = 22444;
	#10 counter$count = 22445;
	#10 counter$count = 22446;
	#10 counter$count = 22447;
	#10 counter$count = 22448;
	#10 counter$count = 22449;
	#10 counter$count = 22450;
	#10 counter$count = 22451;
	#10 counter$count = 22452;
	#10 counter$count = 22453;
	#10 counter$count = 22454;
	#10 counter$count = 22455;
	#10 counter$count = 22456;
	#10 counter$count = 22457;
	#10 counter$count = 22458;
	#10 counter$count = 22459;
	#10 counter$count = 22460;
	#10 counter$count = 22461;
	#10 counter$count = 22462;
	#10 counter$count = 22463;
	#10 counter$count = 22464;
	#10 counter$count = 22465;
	#10 counter$count = 22466;
	#10 counter$count = 22467;
	#10 counter$count = 22468;
	#10 counter$count = 22469;
	#10 counter$count = 22470;
	#10 counter$count = 22471;
	#10 counter$count = 22472;
	#10 counter$count = 22473;
	#10 counter$count = 22474;
	#10 counter$count = 22475;
	#10 counter$count = 22476;
	#10 counter$count = 22477;
	#10 counter$count = 22478;
	#10 counter$count = 22479;
	#10 counter$count = 22480;
	#10 counter$count = 22481;
	#10 counter$count = 22482;
	#10 counter$count = 22483;
	#10 counter$count = 22484;
	#10 counter$count = 22485;
	#10 counter$count = 22486;
	#10 counter$count = 22487;
	#10 counter$count = 22488;
	#10 counter$count = 22489;
	#10 counter$count = 22490;
	#10 counter$count = 22491;
	#10 counter$count = 22492;
	#10 counter$count = 22493;
	#10 counter$count = 22494;
	#10 counter$count = 22495;
	#10 counter$count = 22496;
	#10 counter$count = 22497;
	#10 counter$count = 22498;
	#10 counter$count = 22499;
	#10 counter$count = 22500;
	#10 counter$count = 22501;
	#10 counter$count = 22502;
	#10 counter$count = 22503;
	#10 counter$count = 22504;
	#10 counter$count = 22505;
	#10 counter$count = 22506;
	#10 counter$count = 22507;
	#10 counter$count = 22508;
	#10 counter$count = 22509;
	#10 counter$count = 22510;
	#10 counter$count = 22511;
	#10 counter$count = 22512;
	#10 counter$count = 22513;
	#10 counter$count = 22514;
	#10 counter$count = 22515;
	#10 counter$count = 22516;
	#10 counter$count = 22517;
	#10 counter$count = 22518;
	#10 counter$count = 22519;
	#10 counter$count = 22520;
	#10 counter$count = 22521;
	#10 counter$count = 22522;
	#10 counter$count = 22523;
	#10 counter$count = 22524;
	#10 counter$count = 22525;
	#10 counter$count = 22526;
	#10 counter$count = 22527;
	#10 counter$count = 22528;
	#10 counter$count = 22529;
	#10 counter$count = 22530;
	#10 counter$count = 22531;
	#10 counter$count = 22532;
	#10 counter$count = 22533;
	#10 counter$count = 22534;
	#10 counter$count = 22535;
	#10 counter$count = 22536;
	#10 counter$count = 22537;
	#10 counter$count = 22538;
	#10 counter$count = 22539;
	#10 counter$count = 22540;
	#10 counter$count = 22541;
	#10 counter$count = 22542;
	#10 counter$count = 22543;
	#10 counter$count = 22544;
	#10 counter$count = 22545;
	#10 counter$count = 22546;
	#10 counter$count = 22547;
	#10 counter$count = 22548;
	#10 counter$count = 22549;
	#10 counter$count = 22550;
	#10 counter$count = 22551;
	#10 counter$count = 22552;
	#10 counter$count = 22553;
	#10 counter$count = 22554;
	#10 counter$count = 22555;
	#10 counter$count = 22556;
	#10 counter$count = 22557;
	#10 counter$count = 22558;
	#10 counter$count = 22559;
	#10 counter$count = 22560;
	#10 counter$count = 22561;
	#10 counter$count = 22562;
	#10 counter$count = 22563;
	#10 counter$count = 22564;
	#10 counter$count = 22565;
	#10 counter$count = 22566;
	#10 counter$count = 22567;
	#10 counter$count = 22568;
	#10 counter$count = 22569;
	#10 counter$count = 22570;
	#10 counter$count = 22571;
	#10 counter$count = 22572;
	#10 counter$count = 22573;
	#10 counter$count = 22574;
	#10 counter$count = 22575;
	#10 counter$count = 22576;
	#10 counter$count = 22577;
	#10 counter$count = 22578;
	#10 counter$count = 22579;
	#10 counter$count = 22580;
	#10 counter$count = 22581;
	#10 counter$count = 22582;
	#10 counter$count = 22583;
	#10 counter$count = 22584;
	#10 counter$count = 22585;
	#10 counter$count = 22586;
	#10 counter$count = 22587;
	#10 counter$count = 22588;
	#10 counter$count = 22589;
	#10 counter$count = 22590;
	#10 counter$count = 22591;
	#10 counter$count = 22592;
	#10 counter$count = 22593;
	#10 counter$count = 22594;
	#10 counter$count = 22595;
	#10 counter$count = 22596;
	#10 counter$count = 22597;
	#10 counter$count = 22598;
	#10 counter$count = 22599;
	#10 counter$count = 22600;
	#10 counter$count = 22601;
	#10 counter$count = 22602;
	#10 counter$count = 22603;
	#10 counter$count = 22604;
	#10 counter$count = 22605;
	#10 counter$count = 22606;
	#10 counter$count = 22607;
	#10 counter$count = 22608;
	#10 counter$count = 22609;
	#10 counter$count = 22610;
	#10 counter$count = 22611;
	#10 counter$count = 22612;
	#10 counter$count = 22613;
	#10 counter$count = 22614;
	#10 counter$count = 22615;
	#10 counter$count = 22616;
	#10 counter$count = 22617;
	#10 counter$count = 22618;
	#10 counter$count = 22619;
	#10 counter$count = 22620;
	#10 counter$count = 22621;
	#10 counter$count = 22622;
	#10 counter$count = 22623;
	#10 counter$count = 22624;
	#10 counter$count = 22625;
	#10 counter$count = 22626;
	#10 counter$count = 22627;
	#10 counter$count = 22628;
	#10 counter$count = 22629;
	#10 counter$count = 22630;
	#10 counter$count = 22631;
	#10 counter$count = 22632;
	#10 counter$count = 22633;
	#10 counter$count = 22634;
	#10 counter$count = 22635;
	#10 counter$count = 22636;
	#10 counter$count = 22637;
	#10 counter$count = 22638;
	#10 counter$count = 22639;
	#10 counter$count = 22640;
	#10 counter$count = 22641;
	#10 counter$count = 22642;
	#10 counter$count = 22643;
	#10 counter$count = 22644;
	#10 counter$count = 22645;
	#10 counter$count = 22646;
	#10 counter$count = 22647;
	#10 counter$count = 22648;
	#10 counter$count = 22649;
	#10 counter$count = 22650;
	#10 counter$count = 22651;
	#10 counter$count = 22652;
	#10 counter$count = 22653;
	#10 counter$count = 22654;
	#10 counter$count = 22655;
	#10 counter$count = 22656;
	#10 counter$count = 22657;
	#10 counter$count = 22658;
	#10 counter$count = 22659;
	#10 counter$count = 22660;
	#10 counter$count = 22661;
	#10 counter$count = 22662;
	#10 counter$count = 22663;
	#10 counter$count = 22664;
	#10 counter$count = 22665;
	#10 counter$count = 22666;
	#10 counter$count = 22667;
	#10 counter$count = 22668;
	#10 counter$count = 22669;
	#10 counter$count = 22670;
	#10 counter$count = 22671;
	#10 counter$count = 22672;
	#10 counter$count = 22673;
	#10 counter$count = 22674;
	#10 counter$count = 22675;
	#10 counter$count = 22676;
	#10 counter$count = 22677;
	#10 counter$count = 22678;
	#10 counter$count = 22679;
	#10 counter$count = 22680;
	#10 counter$count = 22681;
	#10 counter$count = 22682;
	#10 counter$count = 22683;
	#10 counter$count = 22684;
	#10 counter$count = 22685;
	#10 counter$count = 22686;
	#10 counter$count = 22687;
	#10 counter$count = 22688;
	#10 counter$count = 22689;
	#10 counter$count = 22690;
	#10 counter$count = 22691;
	#10 counter$count = 22692;
	#10 counter$count = 22693;
	#10 counter$count = 22694;
	#10 counter$count = 22695;
	#10 counter$count = 22696;
	#10 counter$count = 22697;
	#10 counter$count = 22698;
	#10 counter$count = 22699;
	#10 counter$count = 22700;
	#10 counter$count = 22701;
	#10 counter$count = 22702;
	#10 counter$count = 22703;
	#10 counter$count = 22704;
	#10 counter$count = 22705;
	#10 counter$count = 22706;
	#10 counter$count = 22707;
	#10 counter$count = 22708;
	#10 counter$count = 22709;
	#10 counter$count = 22710;
	#10 counter$count = 22711;
	#10 counter$count = 22712;
	#10 counter$count = 22713;
	#10 counter$count = 22714;
	#10 counter$count = 22715;
	#10 counter$count = 22716;
	#10 counter$count = 22717;
	#10 counter$count = 22718;
	#10 counter$count = 22719;
	#10 counter$count = 22720;
	#10 counter$count = 22721;
	#10 counter$count = 22722;
	#10 counter$count = 22723;
	#10 counter$count = 22724;
	#10 counter$count = 22725;
	#10 counter$count = 22726;
	#10 counter$count = 22727;
	#10 counter$count = 22728;
	#10 counter$count = 22729;
	#10 counter$count = 22730;
	#10 counter$count = 22731;
	#10 counter$count = 22732;
	#10 counter$count = 22733;
	#10 counter$count = 22734;
	#10 counter$count = 22735;
	#10 counter$count = 22736;
	#10 counter$count = 22737;
	#10 counter$count = 22738;
	#10 counter$count = 22739;
	#10 counter$count = 22740;
	#10 counter$count = 22741;
	#10 counter$count = 22742;
	#10 counter$count = 22743;
	#10 counter$count = 22744;
	#10 counter$count = 22745;
	#10 counter$count = 22746;
	#10 counter$count = 22747;
	#10 counter$count = 22748;
	#10 counter$count = 22749;
	#10 counter$count = 22750;
	#10 counter$count = 22751;
	#10 counter$count = 22752;
	#10 counter$count = 22753;
	#10 counter$count = 22754;
	#10 counter$count = 22755;
	#10 counter$count = 22756;
	#10 counter$count = 22757;
	#10 counter$count = 22758;
	#10 counter$count = 22759;
	#10 counter$count = 22760;
	#10 counter$count = 22761;
	#10 counter$count = 22762;
	#10 counter$count = 22763;
	#10 counter$count = 22764;
	#10 counter$count = 22765;
	#10 counter$count = 22766;
	#10 counter$count = 22767;
	#10 counter$count = 22768;
	#10 counter$count = 22769;
	#10 counter$count = 22770;
	#10 counter$count = 22771;
	#10 counter$count = 22772;
	#10 counter$count = 22773;
	#10 counter$count = 22774;
	#10 counter$count = 22775;
	#10 counter$count = 22776;
	#10 counter$count = 22777;
	#10 counter$count = 22778;
	#10 counter$count = 22779;
	#10 counter$count = 22780;
	#10 counter$count = 22781;
	#10 counter$count = 22782;
	#10 counter$count = 22783;
	#10 counter$count = 22784;
	#10 counter$count = 22785;
	#10 counter$count = 22786;
	#10 counter$count = 22787;
	#10 counter$count = 22788;
	#10 counter$count = 22789;
	#10 counter$count = 22790;
	#10 counter$count = 22791;
	#10 counter$count = 22792;
	#10 counter$count = 22793;
	#10 counter$count = 22794;
	#10 counter$count = 22795;
	#10 counter$count = 22796;
	#10 counter$count = 22797;
	#10 counter$count = 22798;
	#10 counter$count = 22799;
	#10 counter$count = 22800;
	#10 counter$count = 22801;
	#10 counter$count = 22802;
	#10 counter$count = 22803;
	#10 counter$count = 22804;
	#10 counter$count = 22805;
	#10 counter$count = 22806;
	#10 counter$count = 22807;
	#10 counter$count = 22808;
	#10 counter$count = 22809;
	#10 counter$count = 22810;
	#10 counter$count = 22811;
	#10 counter$count = 22812;
	#10 counter$count = 22813;
	#10 counter$count = 22814;
	#10 counter$count = 22815;
	#10 counter$count = 22816;
	#10 counter$count = 22817;
	#10 counter$count = 22818;
	#10 counter$count = 22819;
	#10 counter$count = 22820;
	#10 counter$count = 22821;
	#10 counter$count = 22822;
	#10 counter$count = 22823;
	#10 counter$count = 22824;
	#10 counter$count = 22825;
	#10 counter$count = 22826;
	#10 counter$count = 22827;
	#10 counter$count = 22828;
	#10 counter$count = 22829;
	#10 counter$count = 22830;
	#10 counter$count = 22831;
	#10 counter$count = 22832;
	#10 counter$count = 22833;
	#10 counter$count = 22834;
	#10 counter$count = 22835;
	#10 counter$count = 22836;
	#10 counter$count = 22837;
	#10 counter$count = 22838;
	#10 counter$count = 22839;
	#10 counter$count = 22840;
	#10 counter$count = 22841;
	#10 counter$count = 22842;
	#10 counter$count = 22843;
	#10 counter$count = 22844;
	#10 counter$count = 22845;
	#10 counter$count = 22846;
	#10 counter$count = 22847;
	#10 counter$count = 22848;
	#10 counter$count = 22849;
	#10 counter$count = 22850;
	#10 counter$count = 22851;
	#10 counter$count = 22852;
	#10 counter$count = 22853;
	#10 counter$count = 22854;
	#10 counter$count = 22855;
	#10 counter$count = 22856;
	#10 counter$count = 22857;
	#10 counter$count = 22858;
	#10 counter$count = 22859;
	#10 counter$count = 22860;
	#10 counter$count = 22861;
	#10 counter$count = 22862;
	#10 counter$count = 22863;
	#10 counter$count = 22864;
	#10 counter$count = 22865;
	#10 counter$count = 22866;
	#10 counter$count = 22867;
	#10 counter$count = 22868;
	#10 counter$count = 22869;
	#10 counter$count = 22870;
	#10 counter$count = 22871;
	#10 counter$count = 22872;
	#10 counter$count = 22873;
	#10 counter$count = 22874;
	#10 counter$count = 22875;
	#10 counter$count = 22876;
	#10 counter$count = 22877;
	#10 counter$count = 22878;
	#10 counter$count = 22879;
	#10 counter$count = 22880;
	#10 counter$count = 22881;
	#10 counter$count = 22882;
	#10 counter$count = 22883;
	#10 counter$count = 22884;
	#10 counter$count = 22885;
	#10 counter$count = 22886;
	#10 counter$count = 22887;
	#10 counter$count = 22888;
	#10 counter$count = 22889;
	#10 counter$count = 22890;
	#10 counter$count = 22891;
	#10 counter$count = 22892;
	#10 counter$count = 22893;
	#10 counter$count = 22894;
	#10 counter$count = 22895;
	#10 counter$count = 22896;
	#10 counter$count = 22897;
	#10 counter$count = 22898;
	#10 counter$count = 22899;
	#10 counter$count = 22900;
	#10 counter$count = 22901;
	#10 counter$count = 22902;
	#10 counter$count = 22903;
	#10 counter$count = 22904;
	#10 counter$count = 22905;
	#10 counter$count = 22906;
	#10 counter$count = 22907;
	#10 counter$count = 22908;
	#10 counter$count = 22909;
	#10 counter$count = 22910;
	#10 counter$count = 22911;
	#10 counter$count = 22912;
	#10 counter$count = 22913;
	#10 counter$count = 22914;
	#10 counter$count = 22915;
	#10 counter$count = 22916;
	#10 counter$count = 22917;
	#10 counter$count = 22918;
	#10 counter$count = 22919;
	#10 counter$count = 22920;
	#10 counter$count = 22921;
	#10 counter$count = 22922;
	#10 counter$count = 22923;
	#10 counter$count = 22924;
	#10 counter$count = 22925;
	#10 counter$count = 22926;
	#10 counter$count = 22927;
	#10 counter$count = 22928;
	#10 counter$count = 22929;
	#10 counter$count = 22930;
	#10 counter$count = 22931;
	#10 counter$count = 22932;
	#10 counter$count = 22933;
	#10 counter$count = 22934;
	#10 counter$count = 22935;
	#10 counter$count = 22936;
	#10 counter$count = 22937;
	#10 counter$count = 22938;
	#10 counter$count = 22939;
	#10 counter$count = 22940;
	#10 counter$count = 22941;
	#10 counter$count = 22942;
	#10 counter$count = 22943;
	#10 counter$count = 22944;
	#10 counter$count = 22945;
	#10 counter$count = 22946;
	#10 counter$count = 22947;
	#10 counter$count = 22948;
	#10 counter$count = 22949;
	#10 counter$count = 22950;
	#10 counter$count = 22951;
	#10 counter$count = 22952;
	#10 counter$count = 22953;
	#10 counter$count = 22954;
	#10 counter$count = 22955;
	#10 counter$count = 22956;
	#10 counter$count = 22957;
	#10 counter$count = 22958;
	#10 counter$count = 22959;
	#10 counter$count = 22960;
	#10 counter$count = 22961;
	#10 counter$count = 22962;
	#10 counter$count = 22963;
	#10 counter$count = 22964;
	#10 counter$count = 22965;
	#10 counter$count = 22966;
	#10 counter$count = 22967;
	#10 counter$count = 22968;
	#10 counter$count = 22969;
	#10 counter$count = 22970;
	#10 counter$count = 22971;
	#10 counter$count = 22972;
	#10 counter$count = 22973;
	#10 counter$count = 22974;
	#10 counter$count = 22975;
	#10 counter$count = 22976;
	#10 counter$count = 22977;
	#10 counter$count = 22978;
	#10 counter$count = 22979;
	#10 counter$count = 22980;
	#10 counter$count = 22981;
	#10 counter$count = 22982;
	#10 counter$count = 22983;
	#10 counter$count = 22984;
	#10 counter$count = 22985;
	#10 counter$count = 22986;
	#10 counter$count = 22987;
	#10 counter$count = 22988;
	#10 counter$count = 22989;
	#10 counter$count = 22990;
	#10 counter$count = 22991;
	#10 counter$count = 22992;
	#10 counter$count = 22993;
	#10 counter$count = 22994;
	#10 counter$count = 22995;
	#10 counter$count = 22996;
	#10 counter$count = 22997;
	#10 counter$count = 22998;
	#10 counter$count = 22999;
	#10 counter$count = 23000;
	#10 counter$count = 23001;
	#10 counter$count = 23002;
	#10 counter$count = 23003;
	#10 counter$count = 23004;
	#10 counter$count = 23005;
	#10 counter$count = 23006;
	#10 counter$count = 23007;
	#10 counter$count = 23008;
	#10 counter$count = 23009;
	#10 counter$count = 23010;
	#10 counter$count = 23011;
	#10 counter$count = 23012;
	#10 counter$count = 23013;
	#10 counter$count = 23014;
	#10 counter$count = 23015;
	#10 counter$count = 23016;
	#10 counter$count = 23017;
	#10 counter$count = 23018;
	#10 counter$count = 23019;
	#10 counter$count = 23020;
	#10 counter$count = 23021;
	#10 counter$count = 23022;
	#10 counter$count = 23023;
	#10 counter$count = 23024;
	#10 counter$count = 23025;
	#10 counter$count = 23026;
	#10 counter$count = 23027;
	#10 counter$count = 23028;
	#10 counter$count = 23029;
	#10 counter$count = 23030;
	#10 counter$count = 23031;
	#10 counter$count = 23032;
	#10 counter$count = 23033;
	#10 counter$count = 23034;
	#10 counter$count = 23035;
	#10 counter$count = 23036;
	#10 counter$count = 23037;
	#10 counter$count = 23038;
	#10 counter$count = 23039;
	#10 counter$count = 23040;
	#10 counter$count = 23041;
	#10 counter$count = 23042;
	#10 counter$count = 23043;
	#10 counter$count = 23044;
	#10 counter$count = 23045;
	#10 counter$count = 23046;
	#10 counter$count = 23047;
	#10 counter$count = 23048;
	#10 counter$count = 23049;
	#10 counter$count = 23050;
	#10 counter$count = 23051;
	#10 counter$count = 23052;
	#10 counter$count = 23053;
	#10 counter$count = 23054;
	#10 counter$count = 23055;
	#10 counter$count = 23056;
	#10 counter$count = 23057;
	#10 counter$count = 23058;
	#10 counter$count = 23059;
	#10 counter$count = 23060;
	#10 counter$count = 23061;
	#10 counter$count = 23062;
	#10 counter$count = 23063;
	#10 counter$count = 23064;
	#10 counter$count = 23065;
	#10 counter$count = 23066;
	#10 counter$count = 23067;
	#10 counter$count = 23068;
	#10 counter$count = 23069;
	#10 counter$count = 23070;
	#10 counter$count = 23071;
	#10 counter$count = 23072;
	#10 counter$count = 23073;
	#10 counter$count = 23074;
	#10 counter$count = 23075;
	#10 counter$count = 23076;
	#10 counter$count = 23077;
	#10 counter$count = 23078;
	#10 counter$count = 23079;
	#10 counter$count = 23080;
	#10 counter$count = 23081;
	#10 counter$count = 23082;
	#10 counter$count = 23083;
	#10 counter$count = 23084;
	#10 counter$count = 23085;
	#10 counter$count = 23086;
	#10 counter$count = 23087;
	#10 counter$count = 23088;
	#10 counter$count = 23089;
	#10 counter$count = 23090;
	#10 counter$count = 23091;
	#10 counter$count = 23092;
	#10 counter$count = 23093;
	#10 counter$count = 23094;
	#10 counter$count = 23095;
	#10 counter$count = 23096;
	#10 counter$count = 23097;
	#10 counter$count = 23098;
	#10 counter$count = 23099;
	#10 counter$count = 23100;
	#10 counter$count = 23101;
	#10 counter$count = 23102;
	#10 counter$count = 23103;
	#10 counter$count = 23104;
	#10 counter$count = 23105;
	#10 counter$count = 23106;
	#10 counter$count = 23107;
	#10 counter$count = 23108;
	#10 counter$count = 23109;
	#10 counter$count = 23110;
	#10 counter$count = 23111;
	#10 counter$count = 23112;
	#10 counter$count = 23113;
	#10 counter$count = 23114;
	#10 counter$count = 23115;
	#10 counter$count = 23116;
	#10 counter$count = 23117;
	#10 counter$count = 23118;
	#10 counter$count = 23119;
	#10 counter$count = 23120;
	#10 counter$count = 23121;
	#10 counter$count = 23122;
	#10 counter$count = 23123;
	#10 counter$count = 23124;
	#10 counter$count = 23125;
	#10 counter$count = 23126;
	#10 counter$count = 23127;
	#10 counter$count = 23128;
	#10 counter$count = 23129;
	#10 counter$count = 23130;
	#10 counter$count = 23131;
	#10 counter$count = 23132;
	#10 counter$count = 23133;
	#10 counter$count = 23134;
	#10 counter$count = 23135;
	#10 counter$count = 23136;
	#10 counter$count = 23137;
	#10 counter$count = 23138;
	#10 counter$count = 23139;
	#10 counter$count = 23140;
	#10 counter$count = 23141;
	#10 counter$count = 23142;
	#10 counter$count = 23143;
	#10 counter$count = 23144;
	#10 counter$count = 23145;
	#10 counter$count = 23146;
	#10 counter$count = 23147;
	#10 counter$count = 23148;
	#10 counter$count = 23149;
	#10 counter$count = 23150;
	#10 counter$count = 23151;
	#10 counter$count = 23152;
	#10 counter$count = 23153;
	#10 counter$count = 23154;
	#10 counter$count = 23155;
	#10 counter$count = 23156;
	#10 counter$count = 23157;
	#10 counter$count = 23158;
	#10 counter$count = 23159;
	#10 counter$count = 23160;
	#10 counter$count = 23161;
	#10 counter$count = 23162;
	#10 counter$count = 23163;
	#10 counter$count = 23164;
	#10 counter$count = 23165;
	#10 counter$count = 23166;
	#10 counter$count = 23167;
	#10 counter$count = 23168;
	#10 counter$count = 23169;
	#10 counter$count = 23170;
	#10 counter$count = 23171;
	#10 counter$count = 23172;
	#10 counter$count = 23173;
	#10 counter$count = 23174;
	#10 counter$count = 23175;
	#10 counter$count = 23176;
	#10 counter$count = 23177;
	#10 counter$count = 23178;
	#10 counter$count = 23179;
	#10 counter$count = 23180;
	#10 counter$count = 23181;
	#10 counter$count = 23182;
	#10 counter$count = 23183;
	#10 counter$count = 23184;
	#10 counter$count = 23185;
	#10 counter$count = 23186;
	#10 counter$count = 23187;
	#10 counter$count = 23188;
	#10 counter$count = 23189;
	#10 counter$count = 23190;
	#10 counter$count = 23191;
	#10 counter$count = 23192;
	#10 counter$count = 23193;
	#10 counter$count = 23194;
	#10 counter$count = 23195;
	#10 counter$count = 23196;
	#10 counter$count = 23197;
	#10 counter$count = 23198;
	#10 counter$count = 23199;
	#10 counter$count = 23200;
	#10 counter$count = 23201;
	#10 counter$count = 23202;
	#10 counter$count = 23203;
	#10 counter$count = 23204;
	#10 counter$count = 23205;
	#10 counter$count = 23206;
	#10 counter$count = 23207;
	#10 counter$count = 23208;
	#10 counter$count = 23209;
	#10 counter$count = 23210;
	#10 counter$count = 23211;
	#10 counter$count = 23212;
	#10 counter$count = 23213;
	#10 counter$count = 23214;
	#10 counter$count = 23215;
	#10 counter$count = 23216;
	#10 counter$count = 23217;
	#10 counter$count = 23218;
	#10 counter$count = 23219;
	#10 counter$count = 23220;
	#10 counter$count = 23221;
	#10 counter$count = 23222;
	#10 counter$count = 23223;
	#10 counter$count = 23224;
	#10 counter$count = 23225;
	#10 counter$count = 23226;
	#10 counter$count = 23227;
	#10 counter$count = 23228;
	#10 counter$count = 23229;
	#10 counter$count = 23230;
	#10 counter$count = 23231;
	#10 counter$count = 23232;
	#10 counter$count = 23233;
	#10 counter$count = 23234;
	#10 counter$count = 23235;
	#10 counter$count = 23236;
	#10 counter$count = 23237;
	#10 counter$count = 23238;
	#10 counter$count = 23239;
	#10 counter$count = 23240;
	#10 counter$count = 23241;
	#10 counter$count = 23242;
	#10 counter$count = 23243;
	#10 counter$count = 23244;
	#10 counter$count = 23245;
	#10 counter$count = 23246;
	#10 counter$count = 23247;
	#10 counter$count = 23248;
	#10 counter$count = 23249;
	#10 counter$count = 23250;
	#10 counter$count = 23251;
	#10 counter$count = 23252;
	#10 counter$count = 23253;
	#10 counter$count = 23254;
	#10 counter$count = 23255;
	#10 counter$count = 23256;
	#10 counter$count = 23257;
	#10 counter$count = 23258;
	#10 counter$count = 23259;
	#10 counter$count = 23260;
	#10 counter$count = 23261;
	#10 counter$count = 23262;
	#10 counter$count = 23263;
	#10 counter$count = 23264;
	#10 counter$count = 23265;
	#10 counter$count = 23266;
	#10 counter$count = 23267;
	#10 counter$count = 23268;
	#10 counter$count = 23269;
	#10 counter$count = 23270;
	#10 counter$count = 23271;
	#10 counter$count = 23272;
	#10 counter$count = 23273;
	#10 counter$count = 23274;
	#10 counter$count = 23275;
	#10 counter$count = 23276;
	#10 counter$count = 23277;
	#10 counter$count = 23278;
	#10 counter$count = 23279;
	#10 counter$count = 23280;
	#10 counter$count = 23281;
	#10 counter$count = 23282;
	#10 counter$count = 23283;
	#10 counter$count = 23284;
	#10 counter$count = 23285;
	#10 counter$count = 23286;
	#10 counter$count = 23287;
	#10 counter$count = 23288;
	#10 counter$count = 23289;
	#10 counter$count = 23290;
	#10 counter$count = 23291;
	#10 counter$count = 23292;
	#10 counter$count = 23293;
	#10 counter$count = 23294;
	#10 counter$count = 23295;
	#10 counter$count = 23296;
	#10 counter$count = 23297;
	#10 counter$count = 23298;
	#10 counter$count = 23299;
	#10 counter$count = 23300;
	#10 counter$count = 23301;
	#10 counter$count = 23302;
	#10 counter$count = 23303;
	#10 counter$count = 23304;
	#10 counter$count = 23305;
	#10 counter$count = 23306;
	#10 counter$count = 23307;
	#10 counter$count = 23308;
	#10 counter$count = 23309;
	#10 counter$count = 23310;
	#10 counter$count = 23311;
	#10 counter$count = 23312;
	#10 counter$count = 23313;
	#10 counter$count = 23314;
	#10 counter$count = 23315;
	#10 counter$count = 23316;
	#10 counter$count = 23317;
	#10 counter$count = 23318;
	#10 counter$count = 23319;
	#10 counter$count = 23320;
	#10 counter$count = 23321;
	#10 counter$count = 23322;
	#10 counter$count = 23323;
	#10 counter$count = 23324;
	#10 counter$count = 23325;
	#10 counter$count = 23326;
	#10 counter$count = 23327;
	#10 counter$count = 23328;
	#10 counter$count = 23329;
	#10 counter$count = 23330;
	#10 counter$count = 23331;
	#10 counter$count = 23332;
	#10 counter$count = 23333;
	#10 counter$count = 23334;
	#10 counter$count = 23335;
	#10 counter$count = 23336;
	#10 counter$count = 23337;
	#10 counter$count = 23338;
	#10 counter$count = 23339;
	#10 counter$count = 23340;
	#10 counter$count = 23341;
	#10 counter$count = 23342;
	#10 counter$count = 23343;
	#10 counter$count = 23344;
	#10 counter$count = 23345;
	#10 counter$count = 23346;
	#10 counter$count = 23347;
	#10 counter$count = 23348;
	#10 counter$count = 23349;
	#10 counter$count = 23350;
	#10 counter$count = 23351;
	#10 counter$count = 23352;
	#10 counter$count = 23353;
	#10 counter$count = 23354;
	#10 counter$count = 23355;
	#10 counter$count = 23356;
	#10 counter$count = 23357;
	#10 counter$count = 23358;
	#10 counter$count = 23359;
	#10 counter$count = 23360;
	#10 counter$count = 23361;
	#10 counter$count = 23362;
	#10 counter$count = 23363;
	#10 counter$count = 23364;
	#10 counter$count = 23365;
	#10 counter$count = 23366;
	#10 counter$count = 23367;
	#10 counter$count = 23368;
	#10 counter$count = 23369;
	#10 counter$count = 23370;
	#10 counter$count = 23371;
	#10 counter$count = 23372;
	#10 counter$count = 23373;
	#10 counter$count = 23374;
	#10 counter$count = 23375;
	#10 counter$count = 23376;
	#10 counter$count = 23377;
	#10 counter$count = 23378;
	#10 counter$count = 23379;
	#10 counter$count = 23380;
	#10 counter$count = 23381;
	#10 counter$count = 23382;
	#10 counter$count = 23383;
	#10 counter$count = 23384;
	#10 counter$count = 23385;
	#10 counter$count = 23386;
	#10 counter$count = 23387;
	#10 counter$count = 23388;
	#10 counter$count = 23389;
	#10 counter$count = 23390;
	#10 counter$count = 23391;
	#10 counter$count = 23392;
	#10 counter$count = 23393;
	#10 counter$count = 23394;
	#10 counter$count = 23395;
	#10 counter$count = 23396;
	#10 counter$count = 23397;
	#10 counter$count = 23398;
	#10 counter$count = 23399;
	#10 counter$count = 23400;
	#10 counter$count = 23401;
	#10 counter$count = 23402;
	#10 counter$count = 23403;
	#10 counter$count = 23404;
	#10 counter$count = 23405;
	#10 counter$count = 23406;
	#10 counter$count = 23407;
	#10 counter$count = 23408;
	#10 counter$count = 23409;
	#10 counter$count = 23410;
	#10 counter$count = 23411;
	#10 counter$count = 23412;
	#10 counter$count = 23413;
	#10 counter$count = 23414;
	#10 counter$count = 23415;
	#10 counter$count = 23416;
	#10 counter$count = 23417;
	#10 counter$count = 23418;
	#10 counter$count = 23419;
	#10 counter$count = 23420;
	#10 counter$count = 23421;
	#10 counter$count = 23422;
	#10 counter$count = 23423;
	#10 counter$count = 23424;
	#10 counter$count = 23425;
	#10 counter$count = 23426;
	#10 counter$count = 23427;
	#10 counter$count = 23428;
	#10 counter$count = 23429;
	#10 counter$count = 23430;
	#10 counter$count = 23431;
	#10 counter$count = 23432;
	#10 counter$count = 23433;
	#10 counter$count = 23434;
	#10 counter$count = 23435;
	#10 counter$count = 23436;
	#10 counter$count = 23437;
	#10 counter$count = 23438;
	#10 counter$count = 23439;
	#10 counter$count = 23440;
	#10 counter$count = 23441;
	#10 counter$count = 23442;
	#10 counter$count = 23443;
	#10 counter$count = 23444;
	#10 counter$count = 23445;
	#10 counter$count = 23446;
	#10 counter$count = 23447;
	#10 counter$count = 23448;
	#10 counter$count = 23449;
	#10 counter$count = 23450;
	#10 counter$count = 23451;
	#10 counter$count = 23452;
	#10 counter$count = 23453;
	#10 counter$count = 23454;
	#10 counter$count = 23455;
	#10 counter$count = 23456;
	#10 counter$count = 23457;
	#10 counter$count = 23458;
	#10 counter$count = 23459;
	#10 counter$count = 23460;
	#10 counter$count = 23461;
	#10 counter$count = 23462;
	#10 counter$count = 23463;
	#10 counter$count = 23464;
	#10 counter$count = 23465;
	#10 counter$count = 23466;
	#10 counter$count = 23467;
	#10 counter$count = 23468;
	#10 counter$count = 23469;
	#10 counter$count = 23470;
	#10 counter$count = 23471;
	#10 counter$count = 23472;
	#10 counter$count = 23473;
	#10 counter$count = 23474;
	#10 counter$count = 23475;
	#10 counter$count = 23476;
	#10 counter$count = 23477;
	#10 counter$count = 23478;
	#10 counter$count = 23479;
	#10 counter$count = 23480;
	#10 counter$count = 23481;
	#10 counter$count = 23482;
	#10 counter$count = 23483;
	#10 counter$count = 23484;
	#10 counter$count = 23485;
	#10 counter$count = 23486;
	#10 counter$count = 23487;
	#10 counter$count = 23488;
	#10 counter$count = 23489;
	#10 counter$count = 23490;
	#10 counter$count = 23491;
	#10 counter$count = 23492;
	#10 counter$count = 23493;
	#10 counter$count = 23494;
	#10 counter$count = 23495;
	#10 counter$count = 23496;
	#10 counter$count = 23497;
	#10 counter$count = 23498;
	#10 counter$count = 23499;
	#10 counter$count = 23500;
	#10 counter$count = 23501;
	#10 counter$count = 23502;
	#10 counter$count = 23503;
	#10 counter$count = 23504;
	#10 counter$count = 23505;
	#10 counter$count = 23506;
	#10 counter$count = 23507;
	#10 counter$count = 23508;
	#10 counter$count = 23509;
	#10 counter$count = 23510;
	#10 counter$count = 23511;
	#10 counter$count = 23512;
	#10 counter$count = 23513;
	#10 counter$count = 23514;
	#10 counter$count = 23515;
	#10 counter$count = 23516;
	#10 counter$count = 23517;
	#10 counter$count = 23518;
	#10 counter$count = 23519;
	#10 counter$count = 23520;
	#10 counter$count = 23521;
	#10 counter$count = 23522;
	#10 counter$count = 23523;
	#10 counter$count = 23524;
	#10 counter$count = 23525;
	#10 counter$count = 23526;
	#10 counter$count = 23527;
	#10 counter$count = 23528;
	#10 counter$count = 23529;
	#10 counter$count = 23530;
	#10 counter$count = 23531;
	#10 counter$count = 23532;
	#10 counter$count = 23533;
	#10 counter$count = 23534;
	#10 counter$count = 23535;
	#10 counter$count = 23536;
	#10 counter$count = 23537;
	#10 counter$count = 23538;
	#10 counter$count = 23539;
	#10 counter$count = 23540;
	#10 counter$count = 23541;
	#10 counter$count = 23542;
	#10 counter$count = 23543;
	#10 counter$count = 23544;
	#10 counter$count = 23545;
	#10 counter$count = 23546;
	#10 counter$count = 23547;
	#10 counter$count = 23548;
	#10 counter$count = 23549;
	#10 counter$count = 23550;
	#10 counter$count = 23551;
	#10 counter$count = 23552;
	#10 counter$count = 23553;
	#10 counter$count = 23554;
	#10 counter$count = 23555;
	#10 counter$count = 23556;
	#10 counter$count = 23557;
	#10 counter$count = 23558;
	#10 counter$count = 23559;
	#10 counter$count = 23560;
	#10 counter$count = 23561;
	#10 counter$count = 23562;
	#10 counter$count = 23563;
	#10 counter$count = 23564;
	#10 counter$count = 23565;
	#10 counter$count = 23566;
	#10 counter$count = 23567;
	#10 counter$count = 23568;
	#10 counter$count = 23569;
	#10 counter$count = 23570;
	#10 counter$count = 23571;
	#10 counter$count = 23572;
	#10 counter$count = 23573;
	#10 counter$count = 23574;
	#10 counter$count = 23575;
	#10 counter$count = 23576;
	#10 counter$count = 23577;
	#10 counter$count = 23578;
	#10 counter$count = 23579;
	#10 counter$count = 23580;
	#10 counter$count = 23581;
	#10 counter$count = 23582;
	#10 counter$count = 23583;
	#10 counter$count = 23584;
	#10 counter$count = 23585;
	#10 counter$count = 23586;
	#10 counter$count = 23587;
	#10 counter$count = 23588;
	#10 counter$count = 23589;
	#10 counter$count = 23590;
	#10 counter$count = 23591;
	#10 counter$count = 23592;
	#10 counter$count = 23593;
	#10 counter$count = 23594;
	#10 counter$count = 23595;
	#10 counter$count = 23596;
	#10 counter$count = 23597;
	#10 counter$count = 23598;
	#10 counter$count = 23599;
	#10 counter$count = 23600;
	#10 counter$count = 23601;
	#10 counter$count = 23602;
	#10 counter$count = 23603;
	#10 counter$count = 23604;
	#10 counter$count = 23605;
	#10 counter$count = 23606;
	#10 counter$count = 23607;
	#10 counter$count = 23608;
	#10 counter$count = 23609;
	#10 counter$count = 23610;
	#10 counter$count = 23611;
	#10 counter$count = 23612;
	#10 counter$count = 23613;
	#10 counter$count = 23614;
	#10 counter$count = 23615;
	#10 counter$count = 23616;
	#10 counter$count = 23617;
	#10 counter$count = 23618;
	#10 counter$count = 23619;
	#10 counter$count = 23620;
	#10 counter$count = 23621;
	#10 counter$count = 23622;
	#10 counter$count = 23623;
	#10 counter$count = 23624;
	#10 counter$count = 23625;
	#10 counter$count = 23626;
	#10 counter$count = 23627;
	#10 counter$count = 23628;
	#10 counter$count = 23629;
	#10 counter$count = 23630;
	#10 counter$count = 23631;
	#10 counter$count = 23632;
	#10 counter$count = 23633;
	#10 counter$count = 23634;
	#10 counter$count = 23635;
	#10 counter$count = 23636;
	#10 counter$count = 23637;
	#10 counter$count = 23638;
	#10 counter$count = 23639;
	#10 counter$count = 23640;
	#10 counter$count = 23641;
	#10 counter$count = 23642;
	#10 counter$count = 23643;
	#10 counter$count = 23644;
	#10 counter$count = 23645;
	#10 counter$count = 23646;
	#10 counter$count = 23647;
	#10 counter$count = 23648;
	#10 counter$count = 23649;
	#10 counter$count = 23650;
	#10 counter$count = 23651;
	#10 counter$count = 23652;
	#10 counter$count = 23653;
	#10 counter$count = 23654;
	#10 counter$count = 23655;
	#10 counter$count = 23656;
	#10 counter$count = 23657;
	#10 counter$count = 23658;
	#10 counter$count = 23659;
	#10 counter$count = 23660;
	#10 counter$count = 23661;
	#10 counter$count = 23662;
	#10 counter$count = 23663;
	#10 counter$count = 23664;
	#10 counter$count = 23665;
	#10 counter$count = 23666;
	#10 counter$count = 23667;
	#10 counter$count = 23668;
	#10 counter$count = 23669;
	#10 counter$count = 23670;
	#10 counter$count = 23671;
	#10 counter$count = 23672;
	#10 counter$count = 23673;
	#10 counter$count = 23674;
	#10 counter$count = 23675;
	#10 counter$count = 23676;
	#10 counter$count = 23677;
	#10 counter$count = 23678;
	#10 counter$count = 23679;
	#10 counter$count = 23680;
	#10 counter$count = 23681;
	#10 counter$count = 23682;
	#10 counter$count = 23683;
	#10 counter$count = 23684;
	#10 counter$count = 23685;
	#10 counter$count = 23686;
	#10 counter$count = 23687;
	#10 counter$count = 23688;
	#10 counter$count = 23689;
	#10 counter$count = 23690;
	#10 counter$count = 23691;
	#10 counter$count = 23692;
	#10 counter$count = 23693;
	#10 counter$count = 23694;
	#10 counter$count = 23695;
	#10 counter$count = 23696;
	#10 counter$count = 23697;
	#10 counter$count = 23698;
	#10 counter$count = 23699;
	#10 counter$count = 23700;
	#10 counter$count = 23701;
	#10 counter$count = 23702;
	#10 counter$count = 23703;
	#10 counter$count = 23704;
	#10 counter$count = 23705;
	#10 counter$count = 23706;
	#10 counter$count = 23707;
	#10 counter$count = 23708;
	#10 counter$count = 23709;
	#10 counter$count = 23710;
	#10 counter$count = 23711;
	#10 counter$count = 23712;
	#10 counter$count = 23713;
	#10 counter$count = 23714;
	#10 counter$count = 23715;
	#10 counter$count = 23716;
	#10 counter$count = 23717;
	#10 counter$count = 23718;
	#10 counter$count = 23719;
	#10 counter$count = 23720;
	#10 counter$count = 23721;
	#10 counter$count = 23722;
	#10 counter$count = 23723;
	#10 counter$count = 23724;
	#10 counter$count = 23725;
	#10 counter$count = 23726;
	#10 counter$count = 23727;
	#10 counter$count = 23728;
	#10 counter$count = 23729;
	#10 counter$count = 23730;
	#10 counter$count = 23731;
	#10 counter$count = 23732;
	#10 counter$count = 23733;
	#10 counter$count = 23734;
	#10 counter$count = 23735;
	#10 counter$count = 23736;
	#10 counter$count = 23737;
	#10 counter$count = 23738;
	#10 counter$count = 23739;
	#10 counter$count = 23740;
	#10 counter$count = 23741;
	#10 counter$count = 23742;
	#10 counter$count = 23743;
	#10 counter$count = 23744;
	#10 counter$count = 23745;
	#10 counter$count = 23746;
	#10 counter$count = 23747;
	#10 counter$count = 23748;
	#10 counter$count = 23749;
	#10 counter$count = 23750;
	#10 counter$count = 23751;
	#10 counter$count = 23752;
	#10 counter$count = 23753;
	#10 counter$count = 23754;
	#10 counter$count = 23755;
	#10 counter$count = 23756;
	#10 counter$count = 23757;
	#10 counter$count = 23758;
	#10 counter$count = 23759;
	#10 counter$count = 23760;
	#10 counter$count = 23761;
	#10 counter$count = 23762;
	#10 counter$count = 23763;
	#10 counter$count = 23764;
	#10 counter$count = 23765;
	#10 counter$count = 23766;
	#10 counter$count = 23767;
	#10 counter$count = 23768;
	#10 counter$count = 23769;
	#10 counter$count = 23770;
	#10 counter$count = 23771;
	#10 counter$count = 23772;
	#10 counter$count = 23773;
	#10 counter$count = 23774;
	#10 counter$count = 23775;
	#10 counter$count = 23776;
	#10 counter$count = 23777;
	#10 counter$count = 23778;
	#10 counter$count = 23779;
	#10 counter$count = 23780;
	#10 counter$count = 23781;
	#10 counter$count = 23782;
	#10 counter$count = 23783;
	#10 counter$count = 23784;
	#10 counter$count = 23785;
	#10 counter$count = 23786;
	#10 counter$count = 23787;
	#10 counter$count = 23788;
	#10 counter$count = 23789;
	#10 counter$count = 23790;
	#10 counter$count = 23791;
	#10 counter$count = 23792;
	#10 counter$count = 23793;
	#10 counter$count = 23794;
	#10 counter$count = 23795;
	#10 counter$count = 23796;
	#10 counter$count = 23797;
	#10 counter$count = 23798;
	#10 counter$count = 23799;
	#10 counter$count = 23800;
	#10 counter$count = 23801;
	#10 counter$count = 23802;
	#10 counter$count = 23803;
	#10 counter$count = 23804;
	#10 counter$count = 23805;
	#10 counter$count = 23806;
	#10 counter$count = 23807;
	#10 counter$count = 23808;
	#10 counter$count = 23809;
	#10 counter$count = 23810;
	#10 counter$count = 23811;
	#10 counter$count = 23812;
	#10 counter$count = 23813;
	#10 counter$count = 23814;
	#10 counter$count = 23815;
	#10 counter$count = 23816;
	#10 counter$count = 23817;
	#10 counter$count = 23818;
	#10 counter$count = 23819;
	#10 counter$count = 23820;
	#10 counter$count = 23821;
	#10 counter$count = 23822;
	#10 counter$count = 23823;
	#10 counter$count = 23824;
	#10 counter$count = 23825;
	#10 counter$count = 23826;
	#10 counter$count = 23827;
	#10 counter$count = 23828;
	#10 counter$count = 23829;
	#10 counter$count = 23830;
	#10 counter$count = 23831;
	#10 counter$count = 23832;
	#10 counter$count = 23833;
	#10 counter$count = 23834;
	#10 counter$count = 23835;
	#10 counter$count = 23836;
	#10 counter$count = 23837;
	#10 counter$count = 23838;
	#10 counter$count = 23839;
	#10 counter$count = 23840;
	#10 counter$count = 23841;
	#10 counter$count = 23842;
	#10 counter$count = 23843;
	#10 counter$count = 23844;
	#10 counter$count = 23845;
	#10 counter$count = 23846;
	#10 counter$count = 23847;
	#10 counter$count = 23848;
	#10 counter$count = 23849;
	#10 counter$count = 23850;
	#10 counter$count = 23851;
	#10 counter$count = 23852;
	#10 counter$count = 23853;
	#10 counter$count = 23854;
	#10 counter$count = 23855;
	#10 counter$count = 23856;
	#10 counter$count = 23857;
	#10 counter$count = 23858;
	#10 counter$count = 23859;
	#10 counter$count = 23860;
	#10 counter$count = 23861;
	#10 counter$count = 23862;
	#10 counter$count = 23863;
	#10 counter$count = 23864;
	#10 counter$count = 23865;
	#10 counter$count = 23866;
	#10 counter$count = 23867;
	#10 counter$count = 23868;
	#10 counter$count = 23869;
	#10 counter$count = 23870;
	#10 counter$count = 23871;
	#10 counter$count = 23872;
	#10 counter$count = 23873;
	#10 counter$count = 23874;
	#10 counter$count = 23875;
	#10 counter$count = 23876;
	#10 counter$count = 23877;
	#10 counter$count = 23878;
	#10 counter$count = 23879;
	#10 counter$count = 23880;
	#10 counter$count = 23881;
	#10 counter$count = 23882;
	#10 counter$count = 23883;
	#10 counter$count = 23884;
	#10 counter$count = 23885;
	#10 counter$count = 23886;
	#10 counter$count = 23887;
	#10 counter$count = 23888;
	#10 counter$count = 23889;
	#10 counter$count = 23890;
	#10 counter$count = 23891;
	#10 counter$count = 23892;
	#10 counter$count = 23893;
	#10 counter$count = 23894;
	#10 counter$count = 23895;
	#10 counter$count = 23896;
	#10 counter$count = 23897;
	#10 counter$count = 23898;
	#10 counter$count = 23899;
	#10 counter$count = 23900;
	#10 counter$count = 23901;
	#10 counter$count = 23902;
	#10 counter$count = 23903;
	#10 counter$count = 23904;
	#10 counter$count = 23905;
	#10 counter$count = 23906;
	#10 counter$count = 23907;
	#10 counter$count = 23908;
	#10 counter$count = 23909;
	#10 counter$count = 23910;
	#10 counter$count = 23911;
	#10 counter$count = 23912;
	#10 counter$count = 23913;
	#10 counter$count = 23914;
	#10 counter$count = 23915;
	#10 counter$count = 23916;
	#10 counter$count = 23917;
	#10 counter$count = 23918;
	#10 counter$count = 23919;
	#10 counter$count = 23920;
	#10 counter$count = 23921;
	#10 counter$count = 23922;
	#10 counter$count = 23923;
	#10 counter$count = 23924;
	#10 counter$count = 23925;
	#10 counter$count = 23926;
	#10 counter$count = 23927;
	#10 counter$count = 23928;
	#10 counter$count = 23929;
	#10 counter$count = 23930;
	#10 counter$count = 23931;
	#10 counter$count = 23932;
	#10 counter$count = 23933;
	#10 counter$count = 23934;
	#10 counter$count = 23935;
	#10 counter$count = 23936;
	#10 counter$count = 23937;
	#10 counter$count = 23938;
	#10 counter$count = 23939;
	#10 counter$count = 23940;
	#10 counter$count = 23941;
	#10 counter$count = 23942;
	#10 counter$count = 23943;
	#10 counter$count = 23944;
	#10 counter$count = 23945;
	#10 counter$count = 23946;
	#10 counter$count = 23947;
	#10 counter$count = 23948;
	#10 counter$count = 23949;
	#10 counter$count = 23950;
	#10 counter$count = 23951;
	#10 counter$count = 23952;
	#10 counter$count = 23953;
	#10 counter$count = 23954;
	#10 counter$count = 23955;
	#10 counter$count = 23956;
	#10 counter$count = 23957;
	#10 counter$count = 23958;
	#10 counter$count = 23959;
	#10 counter$count = 23960;
	#10 counter$count = 23961;
	#10 counter$count = 23962;
	#10 counter$count = 23963;
	#10 counter$count = 23964;
	#10 counter$count = 23965;
	#10 counter$count = 23966;
	#10 counter$count = 23967;
	#10 counter$count = 23968;
	#10 counter$count = 23969;
	#10 counter$count = 23970;
	#10 counter$count = 23971;
	#10 counter$count = 23972;
	#10 counter$count = 23973;
	#10 counter$count = 23974;
	#10 counter$count = 23975;
	#10 counter$count = 23976;
	#10 counter$count = 23977;
	#10 counter$count = 23978;
	#10 counter$count = 23979;
	#10 counter$count = 23980;
	#10 counter$count = 23981;
	#10 counter$count = 23982;
	#10 counter$count = 23983;
	#10 counter$count = 23984;
	#10 counter$count = 23985;
	#10 counter$count = 23986;
	#10 counter$count = 23987;
	#10 counter$count = 23988;
	#10 counter$count = 23989;
	#10 counter$count = 23990;
	#10 counter$count = 23991;
	#10 counter$count = 23992;
	#10 counter$count = 23993;
	#10 counter$count = 23994;
	#10 counter$count = 23995;
	#10 counter$count = 23996;
	#10 counter$count = 23997;
	#10 counter$count = 23998;
	#10 counter$count = 23999;
	#10 counter$count = 24000;
	#10 counter$count = 24001;
	#10 counter$count = 24002;
	#10 counter$count = 24003;
	#10 counter$count = 24004;
	#10 counter$count = 24005;
	#10 counter$count = 24006;
	#10 counter$count = 24007;
	#10 counter$count = 24008;
	#10 counter$count = 24009;
	#10 counter$count = 24010;
	#10 counter$count = 24011;
	#10 counter$count = 24012;
	#10 counter$count = 24013;
	#10 counter$count = 24014;
	#10 counter$count = 24015;
	#10 counter$count = 24016;
	#10 counter$count = 24017;
	#10 counter$count = 24018;
	#10 counter$count = 24019;
	#10 counter$count = 24020;
	#10 counter$count = 24021;
	#10 counter$count = 24022;
	#10 counter$count = 24023;
	#10 counter$count = 24024;
	#10 counter$count = 24025;
	#10 counter$count = 24026;
	#10 counter$count = 24027;
	#10 counter$count = 24028;
	#10 counter$count = 24029;
	#10 counter$count = 24030;
	#10 counter$count = 24031;
	#10 counter$count = 24032;
	#10 counter$count = 24033;
	#10 counter$count = 24034;
	#10 counter$count = 24035;
	#10 counter$count = 24036;
	#10 counter$count = 24037;
	#10 counter$count = 24038;
	#10 counter$count = 24039;
	#10 counter$count = 24040;
	#10 counter$count = 24041;
	#10 counter$count = 24042;
	#10 counter$count = 24043;
	#10 counter$count = 24044;
	#10 counter$count = 24045;
	#10 counter$count = 24046;
	#10 counter$count = 24047;
	#10 counter$count = 24048;
	#10 counter$count = 24049;
	#10 counter$count = 24050;
	#10 counter$count = 24051;
	#10 counter$count = 24052;
	#10 counter$count = 24053;
	#10 counter$count = 24054;
	#10 counter$count = 24055;
	#10 counter$count = 24056;
	#10 counter$count = 24057;
	#10 counter$count = 24058;
	#10 counter$count = 24059;
	#10 counter$count = 24060;
	#10 counter$count = 24061;
	#10 counter$count = 24062;
	#10 counter$count = 24063;
	#10 counter$count = 24064;
	#10 counter$count = 24065;
	#10 counter$count = 24066;
	#10 counter$count = 24067;
	#10 counter$count = 24068;
	#10 counter$count = 24069;
	#10 counter$count = 24070;
	#10 counter$count = 24071;
	#10 counter$count = 24072;
	#10 counter$count = 24073;
	#10 counter$count = 24074;
	#10 counter$count = 24075;
	#10 counter$count = 24076;
	#10 counter$count = 24077;
	#10 counter$count = 24078;
	#10 counter$count = 24079;
	#10 counter$count = 24080;
	#10 counter$count = 24081;
	#10 counter$count = 24082;
	#10 counter$count = 24083;
	#10 counter$count = 24084;
	#10 counter$count = 24085;
	#10 counter$count = 24086;
	#10 counter$count = 24087;
	#10 counter$count = 24088;
	#10 counter$count = 24089;
	#10 counter$count = 24090;
	#10 counter$count = 24091;
	#10 counter$count = 24092;
	#10 counter$count = 24093;
	#10 counter$count = 24094;
	#10 counter$count = 24095;
	#10 counter$count = 24096;
	#10 counter$count = 24097;
	#10 counter$count = 24098;
	#10 counter$count = 24099;
	#10 counter$count = 24100;
	#10 counter$count = 24101;
	#10 counter$count = 24102;
	#10 counter$count = 24103;
	#10 counter$count = 24104;
	#10 counter$count = 24105;
	#10 counter$count = 24106;
	#10 counter$count = 24107;
	#10 counter$count = 24108;
	#10 counter$count = 24109;
	#10 counter$count = 24110;
	#10 counter$count = 24111;
	#10 counter$count = 24112;
	#10 counter$count = 24113;
	#10 counter$count = 24114;
	#10 counter$count = 24115;
	#10 counter$count = 24116;
	#10 counter$count = 24117;
	#10 counter$count = 24118;
	#10 counter$count = 24119;
	#10 counter$count = 24120;
	#10 counter$count = 24121;
	#10 counter$count = 24122;
	#10 counter$count = 24123;
	#10 counter$count = 24124;
	#10 counter$count = 24125;
	#10 counter$count = 24126;
	#10 counter$count = 24127;
	#10 counter$count = 24128;
	#10 counter$count = 24129;
	#10 counter$count = 24130;
	#10 counter$count = 24131;
	#10 counter$count = 24132;
	#10 counter$count = 24133;
	#10 counter$count = 24134;
	#10 counter$count = 24135;
	#10 counter$count = 24136;
	#10 counter$count = 24137;
	#10 counter$count = 24138;
	#10 counter$count = 24139;
	#10 counter$count = 24140;
	#10 counter$count = 24141;
	#10 counter$count = 24142;
	#10 counter$count = 24143;
	#10 counter$count = 24144;
	#10 counter$count = 24145;
	#10 counter$count = 24146;
	#10 counter$count = 24147;
	#10 counter$count = 24148;
	#10 counter$count = 24149;
	#10 counter$count = 24150;
	#10 counter$count = 24151;
	#10 counter$count = 24152;
	#10 counter$count = 24153;
	#10 counter$count = 24154;
	#10 counter$count = 24155;
	#10 counter$count = 24156;
	#10 counter$count = 24157;
	#10 counter$count = 24158;
	#10 counter$count = 24159;
	#10 counter$count = 24160;
	#10 counter$count = 24161;
	#10 counter$count = 24162;
	#10 counter$count = 24163;
	#10 counter$count = 24164;
	#10 counter$count = 24165;
	#10 counter$count = 24166;
	#10 counter$count = 24167;
	#10 counter$count = 24168;
	#10 counter$count = 24169;
	#10 counter$count = 24170;
	#10 counter$count = 24171;
	#10 counter$count = 24172;
	#10 counter$count = 24173;
	#10 counter$count = 24174;
	#10 counter$count = 24175;
	#10 counter$count = 24176;
	#10 counter$count = 24177;
	#10 counter$count = 24178;
	#10 counter$count = 24179;
	#10 counter$count = 24180;
	#10 counter$count = 24181;
	#10 counter$count = 24182;
	#10 counter$count = 24183;
	#10 counter$count = 24184;
	#10 counter$count = 24185;
	#10 counter$count = 24186;
	#10 counter$count = 24187;
	#10 counter$count = 24188;
	#10 counter$count = 24189;
	#10 counter$count = 24190;
	#10 counter$count = 24191;
	#10 counter$count = 24192;
	#10 counter$count = 24193;
	#10 counter$count = 24194;
	#10 counter$count = 24195;
	#10 counter$count = 24196;
	#10 counter$count = 24197;
	#10 counter$count = 24198;
	#10 counter$count = 24199;
	#10 counter$count = 24200;
	#10 counter$count = 24201;
	#10 counter$count = 24202;
	#10 counter$count = 24203;
	#10 counter$count = 24204;
	#10 counter$count = 24205;
	#10 counter$count = 24206;
	#10 counter$count = 24207;
	#10 counter$count = 24208;
	#10 counter$count = 24209;
	#10 counter$count = 24210;
	#10 counter$count = 24211;
	#10 counter$count = 24212;
	#10 counter$count = 24213;
	#10 counter$count = 24214;
	#10 counter$count = 24215;
	#10 counter$count = 24216;
	#10 counter$count = 24217;
	#10 counter$count = 24218;
	#10 counter$count = 24219;
	#10 counter$count = 24220;
	#10 counter$count = 24221;
	#10 counter$count = 24222;
	#10 counter$count = 24223;
	#10 counter$count = 24224;
	#10 counter$count = 24225;
	#10 counter$count = 24226;
	#10 counter$count = 24227;
	#10 counter$count = 24228;
	#10 counter$count = 24229;
	#10 counter$count = 24230;
	#10 counter$count = 24231;
	#10 counter$count = 24232;
	#10 counter$count = 24233;
	#10 counter$count = 24234;
	#10 counter$count = 24235;
	#10 counter$count = 24236;
	#10 counter$count = 24237;
	#10 counter$count = 24238;
	#10 counter$count = 24239;
	#10 counter$count = 24240;
	#10 counter$count = 24241;
	#10 counter$count = 24242;
	#10 counter$count = 24243;
	#10 counter$count = 24244;
	#10 counter$count = 24245;
	#10 counter$count = 24246;
	#10 counter$count = 24247;
	#10 counter$count = 24248;
	#10 counter$count = 24249;
	#10 counter$count = 24250;
	#10 counter$count = 24251;
	#10 counter$count = 24252;
	#10 counter$count = 24253;
	#10 counter$count = 24254;
	#10 counter$count = 24255;
	#10 counter$count = 24256;
	#10 counter$count = 24257;
	#10 counter$count = 24258;
	#10 counter$count = 24259;
	#10 counter$count = 24260;
	#10 counter$count = 24261;
	#10 counter$count = 24262;
	#10 counter$count = 24263;
	#10 counter$count = 24264;
	#10 counter$count = 24265;
	#10 counter$count = 24266;
	#10 counter$count = 24267;
	#10 counter$count = 24268;
	#10 counter$count = 24269;
	#10 counter$count = 24270;
	#10 counter$count = 24271;
	#10 counter$count = 24272;
	#10 counter$count = 24273;
	#10 counter$count = 24274;
	#10 counter$count = 24275;
	#10 counter$count = 24276;
	#10 counter$count = 24277;
	#10 counter$count = 24278;
	#10 counter$count = 24279;
	#10 counter$count = 24280;
	#10 counter$count = 24281;
	#10 counter$count = 24282;
	#10 counter$count = 24283;
	#10 counter$count = 24284;
	#10 counter$count = 24285;
	#10 counter$count = 24286;
	#10 counter$count = 24287;
	#10 counter$count = 24288;
	#10 counter$count = 24289;
	#10 counter$count = 24290;
	#10 counter$count = 24291;
	#10 counter$count = 24292;
	#10 counter$count = 24293;
	#10 counter$count = 24294;
	#10 counter$count = 24295;
	#10 counter$count = 24296;
	#10 counter$count = 24297;
	#10 counter$count = 24298;
	#10 counter$count = 24299;
	#10 counter$count = 24300;
	#10 counter$count = 24301;
	#10 counter$count = 24302;
	#10 counter$count = 24303;
	#10 counter$count = 24304;
	#10 counter$count = 24305;
	#10 counter$count = 24306;
	#10 counter$count = 24307;
	#10 counter$count = 24308;
	#10 counter$count = 24309;
	#10 counter$count = 24310;
	#10 counter$count = 24311;
	#10 counter$count = 24312;
	#10 counter$count = 24313;
	#10 counter$count = 24314;
	#10 counter$count = 24315;
	#10 counter$count = 24316;
	#10 counter$count = 24317;
	#10 counter$count = 24318;
	#10 counter$count = 24319;
	#10 counter$count = 24320;
	#10 counter$count = 24321;
	#10 counter$count = 24322;
	#10 counter$count = 24323;
	#10 counter$count = 24324;
	#10 counter$count = 24325;
	#10 counter$count = 24326;
	#10 counter$count = 24327;
	#10 counter$count = 24328;
	#10 counter$count = 24329;
	#10 counter$count = 24330;
	#10 counter$count = 24331;
	#10 counter$count = 24332;
	#10 counter$count = 24333;
	#10 counter$count = 24334;
	#10 counter$count = 24335;
	#10 counter$count = 24336;
	#10 counter$count = 24337;
	#10 counter$count = 24338;
	#10 counter$count = 24339;
	#10 counter$count = 24340;
	#10 counter$count = 24341;
	#10 counter$count = 24342;
	#10 counter$count = 24343;
	#10 counter$count = 24344;
	#10 counter$count = 24345;
	#10 counter$count = 24346;
	#10 counter$count = 24347;
	#10 counter$count = 24348;
	#10 counter$count = 24349;
	#10 counter$count = 24350;
	#10 counter$count = 24351;
	#10 counter$count = 24352;
	#10 counter$count = 24353;
	#10 counter$count = 24354;
	#10 counter$count = 24355;
	#10 counter$count = 24356;
	#10 counter$count = 24357;
	#10 counter$count = 24358;
	#10 counter$count = 24359;
	#10 counter$count = 24360;
	#10 counter$count = 24361;
	#10 counter$count = 24362;
	#10 counter$count = 24363;
	#10 counter$count = 24364;
	#10 counter$count = 24365;
	#10 counter$count = 24366;
	#10 counter$count = 24367;
	#10 counter$count = 24368;
	#10 counter$count = 24369;
	#10 counter$count = 24370;
	#10 counter$count = 24371;
	#10 counter$count = 24372;
	#10 counter$count = 24373;
	#10 counter$count = 24374;
	#10 counter$count = 24375;
	#10 counter$count = 24376;
	#10 counter$count = 24377;
	#10 counter$count = 24378;
	#10 counter$count = 24379;
	#10 counter$count = 24380;
	#10 counter$count = 24381;
	#10 counter$count = 24382;
	#10 counter$count = 24383;
	#10 counter$count = 24384;
	#10 counter$count = 24385;
	#10 counter$count = 24386;
	#10 counter$count = 24387;
	#10 counter$count = 24388;
	#10 counter$count = 24389;
	#10 counter$count = 24390;
	#10 counter$count = 24391;
	#10 counter$count = 24392;
	#10 counter$count = 24393;
	#10 counter$count = 24394;
	#10 counter$count = 24395;
	#10 counter$count = 24396;
	#10 counter$count = 24397;
	#10 counter$count = 24398;
	#10 counter$count = 24399;
	#10 counter$count = 24400;
	#10 counter$count = 24401;
	#10 counter$count = 24402;
	#10 counter$count = 24403;
	#10 counter$count = 24404;
	#10 counter$count = 24405;
	#10 counter$count = 24406;
	#10 counter$count = 24407;
	#10 counter$count = 24408;
	#10 counter$count = 24409;
	#10 counter$count = 24410;
	#10 counter$count = 24411;
	#10 counter$count = 24412;
	#10 counter$count = 24413;
	#10 counter$count = 24414;
	#10 counter$count = 24415;
	#10 counter$count = 24416;
	#10 counter$count = 24417;
	#10 counter$count = 24418;
	#10 counter$count = 24419;
	#10 counter$count = 24420;
	#10 counter$count = 24421;
	#10 counter$count = 24422;
	#10 counter$count = 24423;
	#10 counter$count = 24424;
	#10 counter$count = 24425;
	#10 counter$count = 24426;
	#10 counter$count = 24427;
	#10 counter$count = 24428;
	#10 counter$count = 24429;
	#10 counter$count = 24430;
	#10 counter$count = 24431;
	#10 counter$count = 24432;
	#10 counter$count = 24433;
	#10 counter$count = 24434;
	#10 counter$count = 24435;
	#10 counter$count = 24436;
	#10 counter$count = 24437;
	#10 counter$count = 24438;
	#10 counter$count = 24439;
	#10 counter$count = 24440;
	#10 counter$count = 24441;
	#10 counter$count = 24442;
	#10 counter$count = 24443;
	#10 counter$count = 24444;
	#10 counter$count = 24445;
	#10 counter$count = 24446;
	#10 counter$count = 24447;
	#10 counter$count = 24448;
	#10 counter$count = 24449;
	#10 counter$count = 24450;
	#10 counter$count = 24451;
	#10 counter$count = 24452;
	#10 counter$count = 24453;
	#10 counter$count = 24454;
	#10 counter$count = 24455;
	#10 counter$count = 24456;
	#10 counter$count = 24457;
	#10 counter$count = 24458;
	#10 counter$count = 24459;
	#10 counter$count = 24460;
	#10 counter$count = 24461;
	#10 counter$count = 24462;
	#10 counter$count = 24463;
	#10 counter$count = 24464;
	#10 counter$count = 24465;
	#10 counter$count = 24466;
	#10 counter$count = 24467;
	#10 counter$count = 24468;
	#10 counter$count = 24469;
	#10 counter$count = 24470;
	#10 counter$count = 24471;
	#10 counter$count = 24472;
	#10 counter$count = 24473;
	#10 counter$count = 24474;
	#10 counter$count = 24475;
	#10 counter$count = 24476;
	#10 counter$count = 24477;
	#10 counter$count = 24478;
	#10 counter$count = 24479;
	#10 counter$count = 24480;
	#10 counter$count = 24481;
	#10 counter$count = 24482;
	#10 counter$count = 24483;
	#10 counter$count = 24484;
	#10 counter$count = 24485;
	#10 counter$count = 24486;
	#10 counter$count = 24487;
	#10 counter$count = 24488;
	#10 counter$count = 24489;
	#10 counter$count = 24490;
	#10 counter$count = 24491;
	#10 counter$count = 24492;
	#10 counter$count = 24493;
	#10 counter$count = 24494;
	#10 counter$count = 24495;
	#10 counter$count = 24496;
	#10 counter$count = 24497;
	#10 counter$count = 24498;
	#10 counter$count = 24499;
	#10 counter$count = 24500;
	#10 counter$count = 24501;
	#10 counter$count = 24502;
	#10 counter$count = 24503;
	#10 counter$count = 24504;
	#10 counter$count = 24505;
	#10 counter$count = 24506;
	#10 counter$count = 24507;
	#10 counter$count = 24508;
	#10 counter$count = 24509;
	#10 counter$count = 24510;
	#10 counter$count = 24511;
	#10 counter$count = 24512;
	#10 counter$count = 24513;
	#10 counter$count = 24514;
	#10 counter$count = 24515;
	#10 counter$count = 24516;
	#10 counter$count = 24517;
	#10 counter$count = 24518;
	#10 counter$count = 24519;
	#10 counter$count = 24520;
	#10 counter$count = 24521;
	#10 counter$count = 24522;
	#10 counter$count = 24523;
	#10 counter$count = 24524;
	#10 counter$count = 24525;
	#10 counter$count = 24526;
	#10 counter$count = 24527;
	#10 counter$count = 24528;
	#10 counter$count = 24529;
	#10 counter$count = 24530;
	#10 counter$count = 24531;
	#10 counter$count = 24532;
	#10 counter$count = 24533;
	#10 counter$count = 24534;
	#10 counter$count = 24535;
	#10 counter$count = 24536;
	#10 counter$count = 24537;
	#10 counter$count = 24538;
	#10 counter$count = 24539;
	#10 counter$count = 24540;
	#10 counter$count = 24541;
	#10 counter$count = 24542;
	#10 counter$count = 24543;
	#10 counter$count = 24544;
	#10 counter$count = 24545;
	#10 counter$count = 24546;
	#10 counter$count = 24547;
	#10 counter$count = 24548;
	#10 counter$count = 24549;
	#10 counter$count = 24550;
	#10 counter$count = 24551;
	#10 counter$count = 24552;
	#10 counter$count = 24553;
	#10 counter$count = 24554;
	#10 counter$count = 24555;
	#10 counter$count = 24556;
	#10 counter$count = 24557;
	#10 counter$count = 24558;
	#10 counter$count = 24559;
	#10 counter$count = 24560;
	#10 counter$count = 24561;
	#10 counter$count = 24562;
	#10 counter$count = 24563;
	#10 counter$count = 24564;
	#10 counter$count = 24565;
	#10 counter$count = 24566;
	#10 counter$count = 24567;
	#10 counter$count = 24568;
	#10 counter$count = 24569;
	#10 counter$count = 24570;
	#10 counter$count = 24571;
	#10 counter$count = 24572;
	#10 counter$count = 24573;
	#10 counter$count = 24574;
	#10 counter$count = 24575;
	#10 counter$count = 24576;
	#10 counter$count = 24577;
	#10 counter$count = 24578;
	#10 counter$count = 24579;
	#10 counter$count = 24580;
	#10 counter$count = 24581;
	#10 counter$count = 24582;
	#10 counter$count = 24583;
	#10 counter$count = 24584;
	#10 counter$count = 24585;
	#10 counter$count = 24586;
	#10 counter$count = 24587;
	#10 counter$count = 24588;
	#10 counter$count = 24589;
	#10 counter$count = 24590;
	#10 counter$count = 24591;
	#10 counter$count = 24592;
	#10 counter$count = 24593;
	#10 counter$count = 24594;
	#10 counter$count = 24595;
	#10 counter$count = 24596;
	#10 counter$count = 24597;
	#10 counter$count = 24598;
	#10 counter$count = 24599;
	#10 counter$count = 24600;
	#10 counter$count = 24601;
	#10 counter$count = 24602;
	#10 counter$count = 24603;
	#10 counter$count = 24604;
	#10 counter$count = 24605;
	#10 counter$count = 24606;
	#10 counter$count = 24607;
	#10 counter$count = 24608;
	#10 counter$count = 24609;
	#10 counter$count = 24610;
	#10 counter$count = 24611;
	#10 counter$count = 24612;
	#10 counter$count = 24613;
	#10 counter$count = 24614;
	#10 counter$count = 24615;
	#10 counter$count = 24616;
	#10 counter$count = 24617;
	#10 counter$count = 24618;
	#10 counter$count = 24619;
	#10 counter$count = 24620;
	#10 counter$count = 24621;
	#10 counter$count = 24622;
	#10 counter$count = 24623;
	#10 counter$count = 24624;
	#10 counter$count = 24625;
	#10 counter$count = 24626;
	#10 counter$count = 24627;
	#10 counter$count = 24628;
	#10 counter$count = 24629;
	#10 counter$count = 24630;
	#10 counter$count = 24631;
	#10 counter$count = 24632;
	#10 counter$count = 24633;
	#10 counter$count = 24634;
	#10 counter$count = 24635;
	#10 counter$count = 24636;
	#10 counter$count = 24637;
	#10 counter$count = 24638;
	#10 counter$count = 24639;
	#10 counter$count = 24640;
	#10 counter$count = 24641;
	#10 counter$count = 24642;
	#10 counter$count = 24643;
	#10 counter$count = 24644;
	#10 counter$count = 24645;
	#10 counter$count = 24646;
	#10 counter$count = 24647;
	#10 counter$count = 24648;
	#10 counter$count = 24649;
	#10 counter$count = 24650;
	#10 counter$count = 24651;
	#10 counter$count = 24652;
	#10 counter$count = 24653;
	#10 counter$count = 24654;
	#10 counter$count = 24655;
	#10 counter$count = 24656;
	#10 counter$count = 24657;
	#10 counter$count = 24658;
	#10 counter$count = 24659;
	#10 counter$count = 24660;
	#10 counter$count = 24661;
	#10 counter$count = 24662;
	#10 counter$count = 24663;
	#10 counter$count = 24664;
	#10 counter$count = 24665;
	#10 counter$count = 24666;
	#10 counter$count = 24667;
	#10 counter$count = 24668;
	#10 counter$count = 24669;
	#10 counter$count = 24670;
	#10 counter$count = 24671;
	#10 counter$count = 24672;
	#10 counter$count = 24673;
	#10 counter$count = 24674;
	#10 counter$count = 24675;
	#10 counter$count = 24676;
	#10 counter$count = 24677;
	#10 counter$count = 24678;
	#10 counter$count = 24679;
	#10 counter$count = 24680;
	#10 counter$count = 24681;
	#10 counter$count = 24682;
	#10 counter$count = 24683;
	#10 counter$count = 24684;
	#10 counter$count = 24685;
	#10 counter$count = 24686;
	#10 counter$count = 24687;
	#10 counter$count = 24688;
	#10 counter$count = 24689;
	#10 counter$count = 24690;
	#10 counter$count = 24691;
	#10 counter$count = 24692;
	#10 counter$count = 24693;
	#10 counter$count = 24694;
	#10 counter$count = 24695;
	#10 counter$count = 24696;
	#10 counter$count = 24697;
	#10 counter$count = 24698;
	#10 counter$count = 24699;
	#10 counter$count = 24700;
	#10 counter$count = 24701;
	#10 counter$count = 24702;
	#10 counter$count = 24703;
	#10 counter$count = 24704;
	#10 counter$count = 24705;
	#10 counter$count = 24706;
	#10 counter$count = 24707;
	#10 counter$count = 24708;
	#10 counter$count = 24709;
	#10 counter$count = 24710;
	#10 counter$count = 24711;
	#10 counter$count = 24712;
	#10 counter$count = 24713;
	#10 counter$count = 24714;
	#10 counter$count = 24715;
	#10 counter$count = 24716;
	#10 counter$count = 24717;
	#10 counter$count = 24718;
	#10 counter$count = 24719;
	#10 counter$count = 24720;
	#10 counter$count = 24721;
	#10 counter$count = 24722;
	#10 counter$count = 24723;
	#10 counter$count = 24724;
	#10 counter$count = 24725;
	#10 counter$count = 24726;
	#10 counter$count = 24727;
	#10 counter$count = 24728;
	#10 counter$count = 24729;
	#10 counter$count = 24730;
	#10 counter$count = 24731;
	#10 counter$count = 24732;
	#10 counter$count = 24733;
	#10 counter$count = 24734;
	#10 counter$count = 24735;
	#10 counter$count = 24736;
	#10 counter$count = 24737;
	#10 counter$count = 24738;
	#10 counter$count = 24739;
	#10 counter$count = 24740;
	#10 counter$count = 24741;
	#10 counter$count = 24742;
	#10 counter$count = 24743;
	#10 counter$count = 24744;
	#10 counter$count = 24745;
	#10 counter$count = 24746;
	#10 counter$count = 24747;
	#10 counter$count = 24748;
	#10 counter$count = 24749;
	#10 counter$count = 24750;
	#10 counter$count = 24751;
	#10 counter$count = 24752;
	#10 counter$count = 24753;
	#10 counter$count = 24754;
	#10 counter$count = 24755;
	#10 counter$count = 24756;
	#10 counter$count = 24757;
	#10 counter$count = 24758;
	#10 counter$count = 24759;
	#10 counter$count = 24760;
	#10 counter$count = 24761;
	#10 counter$count = 24762;
	#10 counter$count = 24763;
	#10 counter$count = 24764;
	#10 counter$count = 24765;
	#10 counter$count = 24766;
	#10 counter$count = 24767;
	#10 counter$count = 24768;
	#10 counter$count = 24769;
	#10 counter$count = 24770;
	#10 counter$count = 24771;
	#10 counter$count = 24772;
	#10 counter$count = 24773;
	#10 counter$count = 24774;
	#10 counter$count = 24775;
	#10 counter$count = 24776;
	#10 counter$count = 24777;
	#10 counter$count = 24778;
	#10 counter$count = 24779;
	#10 counter$count = 24780;
	#10 counter$count = 24781;
	#10 counter$count = 24782;
	#10 counter$count = 24783;
	#10 counter$count = 24784;
	#10 counter$count = 24785;
	#10 counter$count = 24786;
	#10 counter$count = 24787;
	#10 counter$count = 24788;
	#10 counter$count = 24789;
	#10 counter$count = 24790;
	#10 counter$count = 24791;
	#10 counter$count = 24792;
	#10 counter$count = 24793;
	#10 counter$count = 24794;
	#10 counter$count = 24795;
	#10 counter$count = 24796;
	#10 counter$count = 24797;
	#10 counter$count = 24798;
	#10 counter$count = 24799;
	#10 counter$count = 24800;
	#10 counter$count = 24801;
	#10 counter$count = 24802;
	#10 counter$count = 24803;
	#10 counter$count = 24804;
	#10 counter$count = 24805;
	#10 counter$count = 24806;
	#10 counter$count = 24807;
	#10 counter$count = 24808;
	#10 counter$count = 24809;
	#10 counter$count = 24810;
	#10 counter$count = 24811;
	#10 counter$count = 24812;
	#10 counter$count = 24813;
	#10 counter$count = 24814;
	#10 counter$count = 24815;
	#10 counter$count = 24816;
	#10 counter$count = 24817;
	#10 counter$count = 24818;
	#10 counter$count = 24819;
	#10 counter$count = 24820;
	#10 counter$count = 24821;
	#10 counter$count = 24822;
	#10 counter$count = 24823;
	#10 counter$count = 24824;
	#10 counter$count = 24825;
	#10 counter$count = 24826;
	#10 counter$count = 24827;
	#10 counter$count = 24828;
	#10 counter$count = 24829;
	#10 counter$count = 24830;
	#10 counter$count = 24831;
	#10 counter$count = 24832;
	#10 counter$count = 24833;
	#10 counter$count = 24834;
	#10 counter$count = 24835;
	#10 counter$count = 24836;
	#10 counter$count = 24837;
	#10 counter$count = 24838;
	#10 counter$count = 24839;
	#10 counter$count = 24840;
	#10 counter$count = 24841;
	#10 counter$count = 24842;
	#10 counter$count = 24843;
	#10 counter$count = 24844;
	#10 counter$count = 24845;
	#10 counter$count = 24846;
	#10 counter$count = 24847;
	#10 counter$count = 24848;
	#10 counter$count = 24849;
	#10 counter$count = 24850;
	#10 counter$count = 24851;
	#10 counter$count = 24852;
	#10 counter$count = 24853;
	#10 counter$count = 24854;
	#10 counter$count = 24855;
	#10 counter$count = 24856;
	#10 counter$count = 24857;
	#10 counter$count = 24858;
	#10 counter$count = 24859;
	#10 counter$count = 24860;
	#10 counter$count = 24861;
	#10 counter$count = 24862;
	#10 counter$count = 24863;
	#10 counter$count = 24864;
	#10 counter$count = 24865;
	#10 counter$count = 24866;
	#10 counter$count = 24867;
	#10 counter$count = 24868;
	#10 counter$count = 24869;
	#10 counter$count = 24870;
	#10 counter$count = 24871;
	#10 counter$count = 24872;
	#10 counter$count = 24873;
	#10 counter$count = 24874;
	#10 counter$count = 24875;
	#10 counter$count = 24876;
	#10 counter$count = 24877;
	#10 counter$count = 24878;
	#10 counter$count = 24879;
	#10 counter$count = 24880;
	#10 counter$count = 24881;
	#10 counter$count = 24882;
	#10 counter$count = 24883;
	#10 counter$count = 24884;
	#10 counter$count = 24885;
	#10 counter$count = 24886;
	#10 counter$count = 24887;
	#10 counter$count = 24888;
	#10 counter$count = 24889;
	#10 counter$count = 24890;
	#10 counter$count = 24891;
	#10 counter$count = 24892;
	#10 counter$count = 24893;
	#10 counter$count = 24894;
	#10 counter$count = 24895;
	#10 counter$count = 24896;
	#10 counter$count = 24897;
	#10 counter$count = 24898;
	#10 counter$count = 24899;
	#10 counter$count = 24900;
	#10 counter$count = 24901;
	#10 counter$count = 24902;
	#10 counter$count = 24903;
	#10 counter$count = 24904;
	#10 counter$count = 24905;
	#10 counter$count = 24906;
	#10 counter$count = 24907;
	#10 counter$count = 24908;
	#10 counter$count = 24909;
	#10 counter$count = 24910;
	#10 counter$count = 24911;
	#10 counter$count = 24912;
	#10 counter$count = 24913;
	#10 counter$count = 24914;
	#10 counter$count = 24915;
	#10 counter$count = 24916;
	#10 counter$count = 24917;
	#10 counter$count = 24918;
	#10 counter$count = 24919;
	#10 counter$count = 24920;
	#10 counter$count = 24921;
	#10 counter$count = 24922;
	#10 counter$count = 24923;
	#10 counter$count = 24924;
	#10 counter$count = 24925;
	#10 counter$count = 24926;
	#10 counter$count = 24927;
	#10 counter$count = 24928;
	#10 counter$count = 24929;
	#10 counter$count = 24930;
	#10 counter$count = 24931;
	#10 counter$count = 24932;
	#10 counter$count = 24933;
	#10 counter$count = 24934;
	#10 counter$count = 24935;
	#10 counter$count = 24936;
	#10 counter$count = 24937;
	#10 counter$count = 24938;
	#10 counter$count = 24939;
	#10 counter$count = 24940;
	#10 counter$count = 24941;
	#10 counter$count = 24942;
	#10 counter$count = 24943;
	#10 counter$count = 24944;
	#10 counter$count = 24945;
	#10 counter$count = 24946;
	#10 counter$count = 24947;
	#10 counter$count = 24948;
	#10 counter$count = 24949;
	#10 counter$count = 24950;
	#10 counter$count = 24951;
	#10 counter$count = 24952;
	#10 counter$count = 24953;
	#10 counter$count = 24954;
	#10 counter$count = 24955;
	#10 counter$count = 24956;
	#10 counter$count = 24957;
	#10 counter$count = 24958;
	#10 counter$count = 24959;
	#10 counter$count = 24960;
	#10 counter$count = 24961;
	#10 counter$count = 24962;
	#10 counter$count = 24963;
	#10 counter$count = 24964;
	#10 counter$count = 24965;
	#10 counter$count = 24966;
	#10 counter$count = 24967;
	#10 counter$count = 24968;
	#10 counter$count = 24969;
	#10 counter$count = 24970;
	#10 counter$count = 24971;
	#10 counter$count = 24972;
	#10 counter$count = 24973;
	#10 counter$count = 24974;
	#10 counter$count = 24975;
	#10 counter$count = 24976;
	#10 counter$count = 24977;
	#10 counter$count = 24978;
	#10 counter$count = 24979;
	#10 counter$count = 24980;
	#10 counter$count = 24981;
	#10 counter$count = 24982;
	#10 counter$count = 24983;
	#10 counter$count = 24984;
	#10 counter$count = 24985;
	#10 counter$count = 24986;
	#10 counter$count = 24987;
	#10 counter$count = 24988;
	#10 counter$count = 24989;
	#10 counter$count = 24990;
	#10 counter$count = 24991;
	#10 counter$count = 24992;
	#10 counter$count = 24993;
	#10 counter$count = 24994;
	#10 counter$count = 24995;
	#10 counter$count = 24996;
	#10 counter$count = 24997;
	#10 counter$count = 24998;
	#10 counter$count = 24999;
	#10 counter$count = 25000;
	#10 counter$count = 25001;
	#10 counter$count = 25002;
	#10 counter$count = 25003;
	#10 counter$count = 25004;
	#10 counter$count = 25005;
	#10 counter$count = 25006;
	#10 counter$count = 25007;
	#10 counter$count = 25008;
	#10 counter$count = 25009;
	#10 counter$count = 25010;
	#10 counter$count = 25011;
	#10 counter$count = 25012;
	#10 counter$count = 25013;
	#10 counter$count = 25014;
	#10 counter$count = 25015;
	#10 counter$count = 25016;
	#10 counter$count = 25017;
	#10 counter$count = 25018;
	#10 counter$count = 25019;
	#10 counter$count = 25020;
	#10 counter$count = 25021;
	#10 counter$count = 25022;
	#10 counter$count = 25023;
	#10 counter$count = 25024;
	#10 counter$count = 25025;
	#10 counter$count = 25026;
	#10 counter$count = 25027;
	#10 counter$count = 25028;
	#10 counter$count = 25029;
	#10 counter$count = 25030;
	#10 counter$count = 25031;
	#10 counter$count = 25032;
	#10 counter$count = 25033;
	#10 counter$count = 25034;
	#10 counter$count = 25035;
	#10 counter$count = 25036;
	#10 counter$count = 25037;
	#10 counter$count = 25038;
	#10 counter$count = 25039;
	#10 counter$count = 25040;
	#10 counter$count = 25041;
	#10 counter$count = 25042;
	#10 counter$count = 25043;
	#10 counter$count = 25044;
	#10 counter$count = 25045;
	#10 counter$count = 25046;
	#10 counter$count = 25047;
	#10 counter$count = 25048;
	#10 counter$count = 25049;
	#10 counter$count = 25050;
	#10 counter$count = 25051;
	#10 counter$count = 25052;
	#10 counter$count = 25053;
	#10 counter$count = 25054;
	#10 counter$count = 25055;
	#10 counter$count = 25056;
	#10 counter$count = 25057;
	#10 counter$count = 25058;
	#10 counter$count = 25059;
	#10 counter$count = 25060;
	#10 counter$count = 25061;
	#10 counter$count = 25062;
	#10 counter$count = 25063;
	#10 counter$count = 25064;
	#10 counter$count = 25065;
	#10 counter$count = 25066;
	#10 counter$count = 25067;
	#10 counter$count = 25068;
	#10 counter$count = 25069;
	#10 counter$count = 25070;
	#10 counter$count = 25071;
	#10 counter$count = 25072;
	#10 counter$count = 25073;
	#10 counter$count = 25074;
	#10 counter$count = 25075;
	#10 counter$count = 25076;
	#10 counter$count = 25077;
	#10 counter$count = 25078;
	#10 counter$count = 25079;
	#10 counter$count = 25080;
	#10 counter$count = 25081;
	#10 counter$count = 25082;
	#10 counter$count = 25083;
	#10 counter$count = 25084;
	#10 counter$count = 25085;
	#10 counter$count = 25086;
	#10 counter$count = 25087;
	#10 counter$count = 25088;
	#10 counter$count = 25089;
	#10 counter$count = 25090;
	#10 counter$count = 25091;
	#10 counter$count = 25092;
	#10 counter$count = 25093;
	#10 counter$count = 25094;
	#10 counter$count = 25095;
	#10 counter$count = 25096;
	#10 counter$count = 25097;
	#10 counter$count = 25098;
	#10 counter$count = 25099;
	#10 counter$count = 25100;
	#10 counter$count = 25101;
	#10 counter$count = 25102;
	#10 counter$count = 25103;
	#10 counter$count = 25104;
	#10 counter$count = 25105;
	#10 counter$count = 25106;
	#10 counter$count = 25107;
	#10 counter$count = 25108;
	#10 counter$count = 25109;
	#10 counter$count = 25110;
	#10 counter$count = 25111;
	#10 counter$count = 25112;
	#10 counter$count = 25113;
	#10 counter$count = 25114;
	#10 counter$count = 25115;
	#10 counter$count = 25116;
	#10 counter$count = 25117;
	#10 counter$count = 25118;
	#10 counter$count = 25119;
	#10 counter$count = 25120;
	#10 counter$count = 25121;
	#10 counter$count = 25122;
	#10 counter$count = 25123;
	#10 counter$count = 25124;
	#10 counter$count = 25125;
	#10 counter$count = 25126;
	#10 counter$count = 25127;
	#10 counter$count = 25128;
	#10 counter$count = 25129;
	#10 counter$count = 25130;
	#10 counter$count = 25131;
	#10 counter$count = 25132;
	#10 counter$count = 25133;
	#10 counter$count = 25134;
	#10 counter$count = 25135;
	#10 counter$count = 25136;
	#10 counter$count = 25137;
	#10 counter$count = 25138;
	#10 counter$count = 25139;
	#10 counter$count = 25140;
	#10 counter$count = 25141;
	#10 counter$count = 25142;
	#10 counter$count = 25143;
	#10 counter$count = 25144;
	#10 counter$count = 25145;
	#10 counter$count = 25146;
	#10 counter$count = 25147;
	#10 counter$count = 25148;
	#10 counter$count = 25149;
	#10 counter$count = 25150;
	#10 counter$count = 25151;
	#10 counter$count = 25152;
	#10 counter$count = 25153;
	#10 counter$count = 25154;
	#10 counter$count = 25155;
	#10 counter$count = 25156;
	#10 counter$count = 25157;
	#10 counter$count = 25158;
	#10 counter$count = 25159;
	#10 counter$count = 25160;
	#10 counter$count = 25161;
	#10 counter$count = 25162;
	#10 counter$count = 25163;
	#10 counter$count = 25164;
	#10 counter$count = 25165;
	#10 counter$count = 25166;
	#10 counter$count = 25167;
	#10 counter$count = 25168;
	#10 counter$count = 25169;
	#10 counter$count = 25170;
	#10 counter$count = 25171;
	#10 counter$count = 25172;
	#10 counter$count = 25173;
	#10 counter$count = 25174;
	#10 counter$count = 25175;
	#10 counter$count = 25176;
	#10 counter$count = 25177;
	#10 counter$count = 25178;
	#10 counter$count = 25179;
	#10 counter$count = 25180;
	#10 counter$count = 25181;
	#10 counter$count = 25182;
	#10 counter$count = 25183;
	#10 counter$count = 25184;
	#10 counter$count = 25185;
	#10 counter$count = 25186;
	#10 counter$count = 25187;
	#10 counter$count = 25188;
	#10 counter$count = 25189;
	#10 counter$count = 25190;
	#10 counter$count = 25191;
	#10 counter$count = 25192;
	#10 counter$count = 25193;
	#10 counter$count = 25194;
	#10 counter$count = 25195;
	#10 counter$count = 25196;
	#10 counter$count = 25197;
	#10 counter$count = 25198;
	#10 counter$count = 25199;
	#10 counter$count = 25200;
	#10 counter$count = 25201;
	#10 counter$count = 25202;
	#10 counter$count = 25203;
	#10 counter$count = 25204;
	#10 counter$count = 25205;
	#10 counter$count = 25206;
	#10 counter$count = 25207;
	#10 counter$count = 25208;
	#10 counter$count = 25209;
	#10 counter$count = 25210;
	#10 counter$count = 25211;
	#10 counter$count = 25212;
	#10 counter$count = 25213;
	#10 counter$count = 25214;
	#10 counter$count = 25215;
	#10 counter$count = 25216;
	#10 counter$count = 25217;
	#10 counter$count = 25218;
	#10 counter$count = 25219;
	#10 counter$count = 25220;
	#10 counter$count = 25221;
	#10 counter$count = 25222;
	#10 counter$count = 25223;
	#10 counter$count = 25224;
	#10 counter$count = 25225;
	#10 counter$count = 25226;
	#10 counter$count = 25227;
	#10 counter$count = 25228;
	#10 counter$count = 25229;
	#10 counter$count = 25230;
	#10 counter$count = 25231;
	#10 counter$count = 25232;
	#10 counter$count = 25233;
	#10 counter$count = 25234;
	#10 counter$count = 25235;
	#10 counter$count = 25236;
	#10 counter$count = 25237;
	#10 counter$count = 25238;
	#10 counter$count = 25239;
	#10 counter$count = 25240;
	#10 counter$count = 25241;
	#10 counter$count = 25242;
	#10 counter$count = 25243;
	#10 counter$count = 25244;
	#10 counter$count = 25245;
	#10 counter$count = 25246;
	#10 counter$count = 25247;
	#10 counter$count = 25248;
	#10 counter$count = 25249;
	#10 counter$count = 25250;
	#10 counter$count = 25251;
	#10 counter$count = 25252;
	#10 counter$count = 25253;
	#10 counter$count = 25254;
	#10 counter$count = 25255;
	#10 counter$count = 25256;
	#10 counter$count = 25257;
	#10 counter$count = 25258;
	#10 counter$count = 25259;
	#10 counter$count = 25260;
	#10 counter$count = 25261;
	#10 counter$count = 25262;
	#10 counter$count = 25263;
	#10 counter$count = 25264;
	#10 counter$count = 25265;
	#10 counter$count = 25266;
	#10 counter$count = 25267;
	#10 counter$count = 25268;
	#10 counter$count = 25269;
	#10 counter$count = 25270;
	#10 counter$count = 25271;
	#10 counter$count = 25272;
	#10 counter$count = 25273;
	#10 counter$count = 25274;
	#10 counter$count = 25275;
	#10 counter$count = 25276;
	#10 counter$count = 25277;
	#10 counter$count = 25278;
	#10 counter$count = 25279;
	#10 counter$count = 25280;
	#10 counter$count = 25281;
	#10 counter$count = 25282;
	#10 counter$count = 25283;
	#10 counter$count = 25284;
	#10 counter$count = 25285;
	#10 counter$count = 25286;
	#10 counter$count = 25287;
	#10 counter$count = 25288;
	#10 counter$count = 25289;
	#10 counter$count = 25290;
	#10 counter$count = 25291;
	#10 counter$count = 25292;
	#10 counter$count = 25293;
	#10 counter$count = 25294;
	#10 counter$count = 25295;
	#10 counter$count = 25296;
	#10 counter$count = 25297;
	#10 counter$count = 25298;
	#10 counter$count = 25299;
	#10 counter$count = 25300;
	#10 counter$count = 25301;
	#10 counter$count = 25302;
	#10 counter$count = 25303;
	#10 counter$count = 25304;
	#10 counter$count = 25305;
	#10 counter$count = 25306;
	#10 counter$count = 25307;
	#10 counter$count = 25308;
	#10 counter$count = 25309;
	#10 counter$count = 25310;
	#10 counter$count = 25311;
	#10 counter$count = 25312;
	#10 counter$count = 25313;
	#10 counter$count = 25314;
	#10 counter$count = 25315;
	#10 counter$count = 25316;
	#10 counter$count = 25317;
	#10 counter$count = 25318;
	#10 counter$count = 25319;
	#10 counter$count = 25320;
	#10 counter$count = 25321;
	#10 counter$count = 25322;
	#10 counter$count = 25323;
	#10 counter$count = 25324;
	#10 counter$count = 25325;
	#10 counter$count = 25326;
	#10 counter$count = 25327;
	#10 counter$count = 25328;
	#10 counter$count = 25329;
	#10 counter$count = 25330;
	#10 counter$count = 25331;
	#10 counter$count = 25332;
	#10 counter$count = 25333;
	#10 counter$count = 25334;
	#10 counter$count = 25335;
	#10 counter$count = 25336;
	#10 counter$count = 25337;
	#10 counter$count = 25338;
	#10 counter$count = 25339;
	#10 counter$count = 25340;
	#10 counter$count = 25341;
	#10 counter$count = 25342;
	#10 counter$count = 25343;
	#10 counter$count = 25344;
	#10 counter$count = 25345;
	#10 counter$count = 25346;
	#10 counter$count = 25347;
	#10 counter$count = 25348;
	#10 counter$count = 25349;
	#10 counter$count = 25350;
	#10 counter$count = 25351;
	#10 counter$count = 25352;
	#10 counter$count = 25353;
	#10 counter$count = 25354;
	#10 counter$count = 25355;
	#10 counter$count = 25356;
	#10 counter$count = 25357;
	#10 counter$count = 25358;
	#10 counter$count = 25359;
	#10 counter$count = 25360;
	#10 counter$count = 25361;
	#10 counter$count = 25362;
	#10 counter$count = 25363;
	#10 counter$count = 25364;
	#10 counter$count = 25365;
	#10 counter$count = 25366;
	#10 counter$count = 25367;
	#10 counter$count = 25368;
	#10 counter$count = 25369;
	#10 counter$count = 25370;
	#10 counter$count = 25371;
	#10 counter$count = 25372;
	#10 counter$count = 25373;
	#10 counter$count = 25374;
	#10 counter$count = 25375;
	#10 counter$count = 25376;
	#10 counter$count = 25377;
	#10 counter$count = 25378;
	#10 counter$count = 25379;
	#10 counter$count = 25380;
	#10 counter$count = 25381;
	#10 counter$count = 25382;
	#10 counter$count = 25383;
	#10 counter$count = 25384;
	#10 counter$count = 25385;
	#10 counter$count = 25386;
	#10 counter$count = 25387;
	#10 counter$count = 25388;
	#10 counter$count = 25389;
	#10 counter$count = 25390;
	#10 counter$count = 25391;
	#10 counter$count = 25392;
	#10 counter$count = 25393;
	#10 counter$count = 25394;
	#10 counter$count = 25395;
	#10 counter$count = 25396;
	#10 counter$count = 25397;
	#10 counter$count = 25398;
	#10 counter$count = 25399;
	#10 counter$count = 25400;
	#10 counter$count = 25401;
	#10 counter$count = 25402;
	#10 counter$count = 25403;
	#10 counter$count = 25404;
	#10 counter$count = 25405;
	#10 counter$count = 25406;
	#10 counter$count = 25407;
	#10 counter$count = 25408;
	#10 counter$count = 25409;
	#10 counter$count = 25410;
	#10 counter$count = 25411;
	#10 counter$count = 25412;
	#10 counter$count = 25413;
	#10 counter$count = 25414;
	#10 counter$count = 25415;
	#10 counter$count = 25416;
	#10 counter$count = 25417;
	#10 counter$count = 25418;
	#10 counter$count = 25419;
	#10 counter$count = 25420;
	#10 counter$count = 25421;
	#10 counter$count = 25422;
	#10 counter$count = 25423;
	#10 counter$count = 25424;
	#10 counter$count = 25425;
	#10 counter$count = 25426;
	#10 counter$count = 25427;
	#10 counter$count = 25428;
	#10 counter$count = 25429;
	#10 counter$count = 25430;
	#10 counter$count = 25431;
	#10 counter$count = 25432;
	#10 counter$count = 25433;
	#10 counter$count = 25434;
	#10 counter$count = 25435;
	#10 counter$count = 25436;
	#10 counter$count = 25437;
	#10 counter$count = 25438;
	#10 counter$count = 25439;
	#10 counter$count = 25440;
	#10 counter$count = 25441;
	#10 counter$count = 25442;
	#10 counter$count = 25443;
	#10 counter$count = 25444;
	#10 counter$count = 25445;
	#10 counter$count = 25446;
	#10 counter$count = 25447;
	#10 counter$count = 25448;
	#10 counter$count = 25449;
	#10 counter$count = 25450;
	#10 counter$count = 25451;
	#10 counter$count = 25452;
	#10 counter$count = 25453;
	#10 counter$count = 25454;
	#10 counter$count = 25455;
	#10 counter$count = 25456;
	#10 counter$count = 25457;
	#10 counter$count = 25458;
	#10 counter$count = 25459;
	#10 counter$count = 25460;
	#10 counter$count = 25461;
	#10 counter$count = 25462;
	#10 counter$count = 25463;
	#10 counter$count = 25464;
	#10 counter$count = 25465;
	#10 counter$count = 25466;
	#10 counter$count = 25467;
	#10 counter$count = 25468;
	#10 counter$count = 25469;
	#10 counter$count = 25470;
	#10 counter$count = 25471;
	#10 counter$count = 25472;
	#10 counter$count = 25473;
	#10 counter$count = 25474;
	#10 counter$count = 25475;
	#10 counter$count = 25476;
	#10 counter$count = 25477;
	#10 counter$count = 25478;
	#10 counter$count = 25479;
	#10 counter$count = 25480;
	#10 counter$count = 25481;
	#10 counter$count = 25482;
	#10 counter$count = 25483;
	#10 counter$count = 25484;
	#10 counter$count = 25485;
	#10 counter$count = 25486;
	#10 counter$count = 25487;
	#10 counter$count = 25488;
	#10 counter$count = 25489;
	#10 counter$count = 25490;
	#10 counter$count = 25491;
	#10 counter$count = 25492;
	#10 counter$count = 25493;
	#10 counter$count = 25494;
	#10 counter$count = 25495;
	#10 counter$count = 25496;
	#10 counter$count = 25497;
	#10 counter$count = 25498;
	#10 counter$count = 25499;
	#10 counter$count = 25500;
	#10 counter$count = 25501;
	#10 counter$count = 25502;
	#10 counter$count = 25503;
	#10 counter$count = 25504;
	#10 counter$count = 25505;
	#10 counter$count = 25506;
	#10 counter$count = 25507;
	#10 counter$count = 25508;
	#10 counter$count = 25509;
	#10 counter$count = 25510;
	#10 counter$count = 25511;
	#10 counter$count = 25512;
	#10 counter$count = 25513;
	#10 counter$count = 25514;
	#10 counter$count = 25515;
	#10 counter$count = 25516;
	#10 counter$count = 25517;
	#10 counter$count = 25518;
	#10 counter$count = 25519;
	#10 counter$count = 25520;
	#10 counter$count = 25521;
	#10 counter$count = 25522;
	#10 counter$count = 25523;
	#10 counter$count = 25524;
	#10 counter$count = 25525;
	#10 counter$count = 25526;
	#10 counter$count = 25527;
	#10 counter$count = 25528;
	#10 counter$count = 25529;
	#10 counter$count = 25530;
	#10 counter$count = 25531;
	#10 counter$count = 25532;
	#10 counter$count = 25533;
	#10 counter$count = 25534;
	#10 counter$count = 25535;
	#10 counter$count = 25536;
	#10 counter$count = 25537;
	#10 counter$count = 25538;
	#10 counter$count = 25539;
	#10 counter$count = 25540;
	#10 counter$count = 25541;
	#10 counter$count = 25542;
	#10 counter$count = 25543;
	#10 counter$count = 25544;
	#10 counter$count = 25545;
	#10 counter$count = 25546;
	#10 counter$count = 25547;
	#10 counter$count = 25548;
	#10 counter$count = 25549;
	#10 counter$count = 25550;
	#10 counter$count = 25551;
	#10 counter$count = 25552;
	#10 counter$count = 25553;
	#10 counter$count = 25554;
	#10 counter$count = 25555;
	#10 counter$count = 25556;
	#10 counter$count = 25557;
	#10 counter$count = 25558;
	#10 counter$count = 25559;
	#10 counter$count = 25560;
	#10 counter$count = 25561;
	#10 counter$count = 25562;
	#10 counter$count = 25563;
	#10 counter$count = 25564;
	#10 counter$count = 25565;
	#10 counter$count = 25566;
	#10 counter$count = 25567;
	#10 counter$count = 25568;
	#10 counter$count = 25569;
	#10 counter$count = 25570;
	#10 counter$count = 25571;
	#10 counter$count = 25572;
	#10 counter$count = 25573;
	#10 counter$count = 25574;
	#10 counter$count = 25575;
	#10 counter$count = 25576;
	#10 counter$count = 25577;
	#10 counter$count = 25578;
	#10 counter$count = 25579;
	#10 counter$count = 25580;
	#10 counter$count = 25581;
	#10 counter$count = 25582;
	#10 counter$count = 25583;
	#10 counter$count = 25584;
	#10 counter$count = 25585;
	#10 counter$count = 25586;
	#10 counter$count = 25587;
	#10 counter$count = 25588;
	#10 counter$count = 25589;
	#10 counter$count = 25590;
	#10 counter$count = 25591;
	#10 counter$count = 25592;
	#10 counter$count = 25593;
	#10 counter$count = 25594;
	#10 counter$count = 25595;
	#10 counter$count = 25596;
	#10 counter$count = 25597;
	#10 counter$count = 25598;
	#10 counter$count = 25599;
	#10 counter$count = 25600;
	#10 counter$count = 25601;
	#10 counter$count = 25602;
	#10 counter$count = 25603;
	#10 counter$count = 25604;
	#10 counter$count = 25605;
	#10 counter$count = 25606;
	#10 counter$count = 25607;
	#10 counter$count = 25608;
	#10 counter$count = 25609;
	#10 counter$count = 25610;
	#10 counter$count = 25611;
	#10 counter$count = 25612;
	#10 counter$count = 25613;
	#10 counter$count = 25614;
	#10 counter$count = 25615;
	#10 counter$count = 25616;
	#10 counter$count = 25617;
	#10 counter$count = 25618;
	#10 counter$count = 25619;
	#10 counter$count = 25620;
	#10 counter$count = 25621;
	#10 counter$count = 25622;
	#10 counter$count = 25623;
	#10 counter$count = 25624;
	#10 counter$count = 25625;
	#10 counter$count = 25626;
	#10 counter$count = 25627;
	#10 counter$count = 25628;
	#10 counter$count = 25629;
	#10 counter$count = 25630;
	#10 counter$count = 25631;
	#10 counter$count = 25632;
	#10 counter$count = 25633;
	#10 counter$count = 25634;
	#10 counter$count = 25635;
	#10 counter$count = 25636;
	#10 counter$count = 25637;
	#10 counter$count = 25638;
	#10 counter$count = 25639;
	#10 counter$count = 25640;
	#10 counter$count = 25641;
	#10 counter$count = 25642;
	#10 counter$count = 25643;
	#10 counter$count = 25644;
	#10 counter$count = 25645;
	#10 counter$count = 25646;
	#10 counter$count = 25647;
	#10 counter$count = 25648;
	#10 counter$count = 25649;
	#10 counter$count = 25650;
	#10 counter$count = 25651;
	#10 counter$count = 25652;
	#10 counter$count = 25653;
	#10 counter$count = 25654;
	#10 counter$count = 25655;
	#10 counter$count = 25656;
	#10 counter$count = 25657;
	#10 counter$count = 25658;
	#10 counter$count = 25659;
	#10 counter$count = 25660;
	#10 counter$count = 25661;
	#10 counter$count = 25662;
	#10 counter$count = 25663;
	#10 counter$count = 25664;
	#10 counter$count = 25665;
	#10 counter$count = 25666;
	#10 counter$count = 25667;
	#10 counter$count = 25668;
	#10 counter$count = 25669;
	#10 counter$count = 25670;
	#10 counter$count = 25671;
	#10 counter$count = 25672;
	#10 counter$count = 25673;
	#10 counter$count = 25674;
	#10 counter$count = 25675;
	#10 counter$count = 25676;
	#10 counter$count = 25677;
	#10 counter$count = 25678;
	#10 counter$count = 25679;
	#10 counter$count = 25680;
	#10 counter$count = 25681;
	#10 counter$count = 25682;
	#10 counter$count = 25683;
	#10 counter$count = 25684;
	#10 counter$count = 25685;
	#10 counter$count = 25686;
	#10 counter$count = 25687;
	#10 counter$count = 25688;
	#10 counter$count = 25689;
	#10 counter$count = 25690;
	#10 counter$count = 25691;
	#10 counter$count = 25692;
	#10 counter$count = 25693;
	#10 counter$count = 25694;
	#10 counter$count = 25695;
	#10 counter$count = 25696;
	#10 counter$count = 25697;
	#10 counter$count = 25698;
	#10 counter$count = 25699;
	#10 counter$count = 25700;
	#10 counter$count = 25701;
	#10 counter$count = 25702;
	#10 counter$count = 25703;
	#10 counter$count = 25704;
	#10 counter$count = 25705;
	#10 counter$count = 25706;
	#10 counter$count = 25707;
	#10 counter$count = 25708;
	#10 counter$count = 25709;
	#10 counter$count = 25710;
	#10 counter$count = 25711;
	#10 counter$count = 25712;
	#10 counter$count = 25713;
	#10 counter$count = 25714;
	#10 counter$count = 25715;
	#10 counter$count = 25716;
	#10 counter$count = 25717;
	#10 counter$count = 25718;
	#10 counter$count = 25719;
	#10 counter$count = 25720;
	#10 counter$count = 25721;
	#10 counter$count = 25722;
	#10 counter$count = 25723;
	#10 counter$count = 25724;
	#10 counter$count = 25725;
	#10 counter$count = 25726;
	#10 counter$count = 25727;
	#10 counter$count = 25728;
	#10 counter$count = 25729;
	#10 counter$count = 25730;
	#10 counter$count = 25731;
	#10 counter$count = 25732;
	#10 counter$count = 25733;
	#10 counter$count = 25734;
	#10 counter$count = 25735;
	#10 counter$count = 25736;
	#10 counter$count = 25737;
	#10 counter$count = 25738;
	#10 counter$count = 25739;
	#10 counter$count = 25740;
	#10 counter$count = 25741;
	#10 counter$count = 25742;
	#10 counter$count = 25743;
	#10 counter$count = 25744;
	#10 counter$count = 25745;
	#10 counter$count = 25746;
	#10 counter$count = 25747;
	#10 counter$count = 25748;
	#10 counter$count = 25749;
	#10 counter$count = 25750;
	#10 counter$count = 25751;
	#10 counter$count = 25752;
	#10 counter$count = 25753;
	#10 counter$count = 25754;
	#10 counter$count = 25755;
	#10 counter$count = 25756;
	#10 counter$count = 25757;
	#10 counter$count = 25758;
	#10 counter$count = 25759;
	#10 counter$count = 25760;
	#10 counter$count = 25761;
	#10 counter$count = 25762;
	#10 counter$count = 25763;
	#10 counter$count = 25764;
	#10 counter$count = 25765;
	#10 counter$count = 25766;
	#10 counter$count = 25767;
	#10 counter$count = 25768;
	#10 counter$count = 25769;
	#10 counter$count = 25770;
	#10 counter$count = 25771;
	#10 counter$count = 25772;
	#10 counter$count = 25773;
	#10 counter$count = 25774;
	#10 counter$count = 25775;
	#10 counter$count = 25776;
	#10 counter$count = 25777;
	#10 counter$count = 25778;
	#10 counter$count = 25779;
	#10 counter$count = 25780;
	#10 counter$count = 25781;
	#10 counter$count = 25782;
	#10 counter$count = 25783;
	#10 counter$count = 25784;
	#10 counter$count = 25785;
	#10 counter$count = 25786;
	#10 counter$count = 25787;
	#10 counter$count = 25788;
	#10 counter$count = 25789;
	#10 counter$count = 25790;
	#10 counter$count = 25791;
	#10 counter$count = 25792;
	#10 counter$count = 25793;
	#10 counter$count = 25794;
	#10 counter$count = 25795;
	#10 counter$count = 25796;
	#10 counter$count = 25797;
	#10 counter$count = 25798;
	#10 counter$count = 25799;
	#10 counter$count = 25800;
	#10 counter$count = 25801;
	#10 counter$count = 25802;
	#10 counter$count = 25803;
	#10 counter$count = 25804;
	#10 counter$count = 25805;
	#10 counter$count = 25806;
	#10 counter$count = 25807;
	#10 counter$count = 25808;
	#10 counter$count = 25809;
	#10 counter$count = 25810;
	#10 counter$count = 25811;
	#10 counter$count = 25812;
	#10 counter$count = 25813;
	#10 counter$count = 25814;
	#10 counter$count = 25815;
	#10 counter$count = 25816;
	#10 counter$count = 25817;
	#10 counter$count = 25818;
	#10 counter$count = 25819;
	#10 counter$count = 25820;
	#10 counter$count = 25821;
	#10 counter$count = 25822;
	#10 counter$count = 25823;
	#10 counter$count = 25824;
	#10 counter$count = 25825;
	#10 counter$count = 25826;
	#10 counter$count = 25827;
	#10 counter$count = 25828;
	#10 counter$count = 25829;
	#10 counter$count = 25830;
	#10 counter$count = 25831;
	#10 counter$count = 25832;
	#10 counter$count = 25833;
	#10 counter$count = 25834;
	#10 counter$count = 25835;
	#10 counter$count = 25836;
	#10 counter$count = 25837;
	#10 counter$count = 25838;
	#10 counter$count = 25839;
	#10 counter$count = 25840;
	#10 counter$count = 25841;
	#10 counter$count = 25842;
	#10 counter$count = 25843;
	#10 counter$count = 25844;
	#10 counter$count = 25845;
	#10 counter$count = 25846;
	#10 counter$count = 25847;
	#10 counter$count = 25848;
	#10 counter$count = 25849;
	#10 counter$count = 25850;
	#10 counter$count = 25851;
	#10 counter$count = 25852;
	#10 counter$count = 25853;
	#10 counter$count = 25854;
	#10 counter$count = 25855;
	#10 counter$count = 25856;
	#10 counter$count = 25857;
	#10 counter$count = 25858;
	#10 counter$count = 25859;
	#10 counter$count = 25860;
	#10 counter$count = 25861;
	#10 counter$count = 25862;
	#10 counter$count = 25863;
	#10 counter$count = 25864;
	#10 counter$count = 25865;
	#10 counter$count = 25866;
	#10 counter$count = 25867;
	#10 counter$count = 25868;
	#10 counter$count = 25869;
	#10 counter$count = 25870;
	#10 counter$count = 25871;
	#10 counter$count = 25872;
	#10 counter$count = 25873;
	#10 counter$count = 25874;
	#10 counter$count = 25875;
	#10 counter$count = 25876;
	#10 counter$count = 25877;
	#10 counter$count = 25878;
	#10 counter$count = 25879;
	#10 counter$count = 25880;
	#10 counter$count = 25881;
	#10 counter$count = 25882;
	#10 counter$count = 25883;
	#10 counter$count = 25884;
	#10 counter$count = 25885;
	#10 counter$count = 25886;
	#10 counter$count = 25887;
	#10 counter$count = 25888;
	#10 counter$count = 25889;
	#10 counter$count = 25890;
	#10 counter$count = 25891;
	#10 counter$count = 25892;
	#10 counter$count = 25893;
	#10 counter$count = 25894;
	#10 counter$count = 25895;
	#10 counter$count = 25896;
	#10 counter$count = 25897;
	#10 counter$count = 25898;
	#10 counter$count = 25899;
	#10 counter$count = 25900;
	#10 counter$count = 25901;
	#10 counter$count = 25902;
	#10 counter$count = 25903;
	#10 counter$count = 25904;
	#10 counter$count = 25905;
	#10 counter$count = 25906;
	#10 counter$count = 25907;
	#10 counter$count = 25908;
	#10 counter$count = 25909;
	#10 counter$count = 25910;
	#10 counter$count = 25911;
	#10 counter$count = 25912;
	#10 counter$count = 25913;
	#10 counter$count = 25914;
	#10 counter$count = 25915;
	#10 counter$count = 25916;
	#10 counter$count = 25917;
	#10 counter$count = 25918;
	#10 counter$count = 25919;
	#10 counter$count = 25920;
	#10 counter$count = 25921;
	#10 counter$count = 25922;
	#10 counter$count = 25923;
	#10 counter$count = 25924;
	#10 counter$count = 25925;
	#10 counter$count = 25926;
	#10 counter$count = 25927;
	#10 counter$count = 25928;
	#10 counter$count = 25929;
	#10 counter$count = 25930;
	#10 counter$count = 25931;
	#10 counter$count = 25932;
	#10 counter$count = 25933;
	#10 counter$count = 25934;
	#10 counter$count = 25935;
	#10 counter$count = 25936;
	#10 counter$count = 25937;
	#10 counter$count = 25938;
	#10 counter$count = 25939;
	#10 counter$count = 25940;
	#10 counter$count = 25941;
	#10 counter$count = 25942;
	#10 counter$count = 25943;
	#10 counter$count = 25944;
	#10 counter$count = 25945;
	#10 counter$count = 25946;
	#10 counter$count = 25947;
	#10 counter$count = 25948;
	#10 counter$count = 25949;
	#10 counter$count = 25950;
	#10 counter$count = 25951;
	#10 counter$count = 25952;
	#10 counter$count = 25953;
	#10 counter$count = 25954;
	#10 counter$count = 25955;
	#10 counter$count = 25956;
	#10 counter$count = 25957;
	#10 counter$count = 25958;
	#10 counter$count = 25959;
	#10 counter$count = 25960;
	#10 counter$count = 25961;
	#10 counter$count = 25962;
	#10 counter$count = 25963;
	#10 counter$count = 25964;
	#10 counter$count = 25965;
	#10 counter$count = 25966;
	#10 counter$count = 25967;
	#10 counter$count = 25968;
	#10 counter$count = 25969;
	#10 counter$count = 25970;
	#10 counter$count = 25971;
	#10 counter$count = 25972;
	#10 counter$count = 25973;
	#10 counter$count = 25974;
	#10 counter$count = 25975;
	#10 counter$count = 25976;
	#10 counter$count = 25977;
	#10 counter$count = 25978;
	#10 counter$count = 25979;
	#10 counter$count = 25980;
	#10 counter$count = 25981;
	#10 counter$count = 25982;
	#10 counter$count = 25983;
	#10 counter$count = 25984;
	#10 counter$count = 25985;
	#10 counter$count = 25986;
	#10 counter$count = 25987;
	#10 counter$count = 25988;
	#10 counter$count = 25989;
	#10 counter$count = 25990;
	#10 counter$count = 25991;
	#10 counter$count = 25992;
	#10 counter$count = 25993;
	#10 counter$count = 25994;
	#10 counter$count = 25995;
	#10 counter$count = 25996;
	#10 counter$count = 25997;
	#10 counter$count = 25998;
	#10 counter$count = 25999;
	#10 counter$count = 26000;
	#10 counter$count = 26001;
	#10 counter$count = 26002;
	#10 counter$count = 26003;
	#10 counter$count = 26004;
	#10 counter$count = 26005;
	#10 counter$count = 26006;
	#10 counter$count = 26007;
	#10 counter$count = 26008;
	#10 counter$count = 26009;
	#10 counter$count = 26010;
	#10 counter$count = 26011;
	#10 counter$count = 26012;
	#10 counter$count = 26013;
	#10 counter$count = 26014;
	#10 counter$count = 26015;
	#10 counter$count = 26016;
	#10 counter$count = 26017;
	#10 counter$count = 26018;
	#10 counter$count = 26019;
	#10 counter$count = 26020;
	#10 counter$count = 26021;
	#10 counter$count = 26022;
	#10 counter$count = 26023;
	#10 counter$count = 26024;
	#10 counter$count = 26025;
	#10 counter$count = 26026;
	#10 counter$count = 26027;
	#10 counter$count = 26028;
	#10 counter$count = 26029;
	#10 counter$count = 26030;
	#10 counter$count = 26031;
	#10 counter$count = 26032;
	#10 counter$count = 26033;
	#10 counter$count = 26034;
	#10 counter$count = 26035;
	#10 counter$count = 26036;
	#10 counter$count = 26037;
	#10 counter$count = 26038;
	#10 counter$count = 26039;
	#10 counter$count = 26040;
	#10 counter$count = 26041;
	#10 counter$count = 26042;
	#10 counter$count = 26043;
	#10 counter$count = 26044;
	#10 counter$count = 26045;
	#10 counter$count = 26046;
	#10 counter$count = 26047;
	#10 counter$count = 26048;
	#10 counter$count = 26049;
	#10 counter$count = 26050;
	#10 counter$count = 26051;
	#10 counter$count = 26052;
	#10 counter$count = 26053;
	#10 counter$count = 26054;
	#10 counter$count = 26055;
	#10 counter$count = 26056;
	#10 counter$count = 26057;
	#10 counter$count = 26058;
	#10 counter$count = 26059;
	#10 counter$count = 26060;
	#10 counter$count = 26061;
	#10 counter$count = 26062;
	#10 counter$count = 26063;
	#10 counter$count = 26064;
	#10 counter$count = 26065;
	#10 counter$count = 26066;
	#10 counter$count = 26067;
	#10 counter$count = 26068;
	#10 counter$count = 26069;
	#10 counter$count = 26070;
	#10 counter$count = 26071;
	#10 counter$count = 26072;
	#10 counter$count = 26073;
	#10 counter$count = 26074;
	#10 counter$count = 26075;
	#10 counter$count = 26076;
	#10 counter$count = 26077;
	#10 counter$count = 26078;
	#10 counter$count = 26079;
	#10 counter$count = 26080;
	#10 counter$count = 26081;
	#10 counter$count = 26082;
	#10 counter$count = 26083;
	#10 counter$count = 26084;
	#10 counter$count = 26085;
	#10 counter$count = 26086;
	#10 counter$count = 26087;
	#10 counter$count = 26088;
	#10 counter$count = 26089;
	#10 counter$count = 26090;
	#10 counter$count = 26091;
	#10 counter$count = 26092;
	#10 counter$count = 26093;
	#10 counter$count = 26094;
	#10 counter$count = 26095;
	#10 counter$count = 26096;
	#10 counter$count = 26097;
	#10 counter$count = 26098;
	#10 counter$count = 26099;
	#10 counter$count = 26100;
	#10 counter$count = 26101;
	#10 counter$count = 26102;
	#10 counter$count = 26103;
	#10 counter$count = 26104;
	#10 counter$count = 26105;
	#10 counter$count = 26106;
	#10 counter$count = 26107;
	#10 counter$count = 26108;
	#10 counter$count = 26109;
	#10 counter$count = 26110;
	#10 counter$count = 26111;
	#10 counter$count = 26112;
	#10 counter$count = 26113;
	#10 counter$count = 26114;
	#10 counter$count = 26115;
	#10 counter$count = 26116;
	#10 counter$count = 26117;
	#10 counter$count = 26118;
	#10 counter$count = 26119;
	#10 counter$count = 26120;
	#10 counter$count = 26121;
	#10 counter$count = 26122;
	#10 counter$count = 26123;
	#10 counter$count = 26124;
	#10 counter$count = 26125;
	#10 counter$count = 26126;
	#10 counter$count = 26127;
	#10 counter$count = 26128;
	#10 counter$count = 26129;
	#10 counter$count = 26130;
	#10 counter$count = 26131;
	#10 counter$count = 26132;
	#10 counter$count = 26133;
	#10 counter$count = 26134;
	#10 counter$count = 26135;
	#10 counter$count = 26136;
	#10 counter$count = 26137;
	#10 counter$count = 26138;
	#10 counter$count = 26139;
	#10 counter$count = 26140;
	#10 counter$count = 26141;
	#10 counter$count = 26142;
	#10 counter$count = 26143;
	#10 counter$count = 26144;
	#10 counter$count = 26145;
	#10 counter$count = 26146;
	#10 counter$count = 26147;
	#10 counter$count = 26148;
	#10 counter$count = 26149;
	#10 counter$count = 26150;
	#10 counter$count = 26151;
	#10 counter$count = 26152;
	#10 counter$count = 26153;
	#10 counter$count = 26154;
	#10 counter$count = 26155;
	#10 counter$count = 26156;
	#10 counter$count = 26157;
	#10 counter$count = 26158;
	#10 counter$count = 26159;
	#10 counter$count = 26160;
	#10 counter$count = 26161;
	#10 counter$count = 26162;
	#10 counter$count = 26163;
	#10 counter$count = 26164;
	#10 counter$count = 26165;
	#10 counter$count = 26166;
	#10 counter$count = 26167;
	#10 counter$count = 26168;
	#10 counter$count = 26169;
	#10 counter$count = 26170;
	#10 counter$count = 26171;
	#10 counter$count = 26172;
	#10 counter$count = 26173;
	#10 counter$count = 26174;
	#10 counter$count = 26175;
	#10 counter$count = 26176;
	#10 counter$count = 26177;
	#10 counter$count = 26178;
	#10 counter$count = 26179;
	#10 counter$count = 26180;
	#10 counter$count = 26181;
	#10 counter$count = 26182;
	#10 counter$count = 26183;
	#10 counter$count = 26184;
	#10 counter$count = 26185;
	#10 counter$count = 26186;
	#10 counter$count = 26187;
	#10 counter$count = 26188;
	#10 counter$count = 26189;
	#10 counter$count = 26190;
	#10 counter$count = 26191;
	#10 counter$count = 26192;
	#10 counter$count = 26193;
	#10 counter$count = 26194;
	#10 counter$count = 26195;
	#10 counter$count = 26196;
	#10 counter$count = 26197;
	#10 counter$count = 26198;
	#10 counter$count = 26199;
	#10 counter$count = 26200;
	#10 counter$count = 26201;
	#10 counter$count = 26202;
	#10 counter$count = 26203;
	#10 counter$count = 26204;
	#10 counter$count = 26205;
	#10 counter$count = 26206;
	#10 counter$count = 26207;
	#10 counter$count = 26208;
	#10 counter$count = 26209;
	#10 counter$count = 26210;
	#10 counter$count = 26211;
	#10 counter$count = 26212;
	#10 counter$count = 26213;
	#10 counter$count = 26214;
	#10 counter$count = 26215;
	#10 counter$count = 26216;
	#10 counter$count = 26217;
	#10 counter$count = 26218;
	#10 counter$count = 26219;
	#10 counter$count = 26220;
	#10 counter$count = 26221;
	#10 counter$count = 26222;
	#10 counter$count = 26223;
	#10 counter$count = 26224;
	#10 counter$count = 26225;
	#10 counter$count = 26226;
	#10 counter$count = 26227;
	#10 counter$count = 26228;
	#10 counter$count = 26229;
	#10 counter$count = 26230;
	#10 counter$count = 26231;
	#10 counter$count = 26232;
	#10 counter$count = 26233;
	#10 counter$count = 26234;
	#10 counter$count = 26235;
	#10 counter$count = 26236;
	#10 counter$count = 26237;
	#10 counter$count = 26238;
	#10 counter$count = 26239;
	#10 counter$count = 26240;
	#10 counter$count = 26241;
	#10 counter$count = 26242;
	#10 counter$count = 26243;
	#10 counter$count = 26244;
	#10 counter$count = 26245;
	#10 counter$count = 26246;
	#10 counter$count = 26247;
	#10 counter$count = 26248;
	#10 counter$count = 26249;
	#10 counter$count = 26250;
	#10 counter$count = 26251;
	#10 counter$count = 26252;
	#10 counter$count = 26253;
	#10 counter$count = 26254;
	#10 counter$count = 26255;
	#10 counter$count = 26256;
	#10 counter$count = 26257;
	#10 counter$count = 26258;
	#10 counter$count = 26259;
	#10 counter$count = 26260;
	#10 counter$count = 26261;
	#10 counter$count = 26262;
	#10 counter$count = 26263;
	#10 counter$count = 26264;
	#10 counter$count = 26265;
	#10 counter$count = 26266;
	#10 counter$count = 26267;
	#10 counter$count = 26268;
	#10 counter$count = 26269;
	#10 counter$count = 26270;
	#10 counter$count = 26271;
	#10 counter$count = 26272;
	#10 counter$count = 26273;
	#10 counter$count = 26274;
	#10 counter$count = 26275;
	#10 counter$count = 26276;
	#10 counter$count = 26277;
	#10 counter$count = 26278;
	#10 counter$count = 26279;
	#10 counter$count = 26280;
	#10 counter$count = 26281;
	#10 counter$count = 26282;
	#10 counter$count = 26283;
	#10 counter$count = 26284;
	#10 counter$count = 26285;
	#10 counter$count = 26286;
	#10 counter$count = 26287;
	#10 counter$count = 26288;
	#10 counter$count = 26289;
	#10 counter$count = 26290;
	#10 counter$count = 26291;
	#10 counter$count = 26292;
	#10 counter$count = 26293;
	#10 counter$count = 26294;
	#10 counter$count = 26295;
	#10 counter$count = 26296;
	#10 counter$count = 26297;
	#10 counter$count = 26298;
	#10 counter$count = 26299;
	#10 counter$count = 26300;
	#10 counter$count = 26301;
	#10 counter$count = 26302;
	#10 counter$count = 26303;
	#10 counter$count = 26304;
	#10 counter$count = 26305;
	#10 counter$count = 26306;
	#10 counter$count = 26307;
	#10 counter$count = 26308;
	#10 counter$count = 26309;
	#10 counter$count = 26310;
	#10 counter$count = 26311;
	#10 counter$count = 26312;
	#10 counter$count = 26313;
	#10 counter$count = 26314;
	#10 counter$count = 26315;
	#10 counter$count = 26316;
	#10 counter$count = 26317;
	#10 counter$count = 26318;
	#10 counter$count = 26319;
	#10 counter$count = 26320;
	#10 counter$count = 26321;
	#10 counter$count = 26322;
	#10 counter$count = 26323;
	#10 counter$count = 26324;
	#10 counter$count = 26325;
	#10 counter$count = 26326;
	#10 counter$count = 26327;
	#10 counter$count = 26328;
	#10 counter$count = 26329;
	#10 counter$count = 26330;
	#10 counter$count = 26331;
	#10 counter$count = 26332;
	#10 counter$count = 26333;
	#10 counter$count = 26334;
	#10 counter$count = 26335;
	#10 counter$count = 26336;
	#10 counter$count = 26337;
	#10 counter$count = 26338;
	#10 counter$count = 26339;
	#10 counter$count = 26340;
	#10 counter$count = 26341;
	#10 counter$count = 26342;
	#10 counter$count = 26343;
	#10 counter$count = 26344;
	#10 counter$count = 26345;
	#10 counter$count = 26346;
	#10 counter$count = 26347;
	#10 counter$count = 26348;
	#10 counter$count = 26349;
	#10 counter$count = 26350;
	#10 counter$count = 26351;
	#10 counter$count = 26352;
	#10 counter$count = 26353;
	#10 counter$count = 26354;
	#10 counter$count = 26355;
	#10 counter$count = 26356;
	#10 counter$count = 26357;
	#10 counter$count = 26358;
	#10 counter$count = 26359;
	#10 counter$count = 26360;
	#10 counter$count = 26361;
	#10 counter$count = 26362;
	#10 counter$count = 26363;
	#10 counter$count = 26364;
	#10 counter$count = 26365;
	#10 counter$count = 26366;
	#10 counter$count = 26367;
	#10 counter$count = 26368;
	#10 counter$count = 26369;
	#10 counter$count = 26370;
	#10 counter$count = 26371;
	#10 counter$count = 26372;
	#10 counter$count = 26373;
	#10 counter$count = 26374;
	#10 counter$count = 26375;
	#10 counter$count = 26376;
	#10 counter$count = 26377;
	#10 counter$count = 26378;
	#10 counter$count = 26379;
	#10 counter$count = 26380;
	#10 counter$count = 26381;
	#10 counter$count = 26382;
	#10 counter$count = 26383;
	#10 counter$count = 26384;
	#10 counter$count = 26385;
	#10 counter$count = 26386;
	#10 counter$count = 26387;
	#10 counter$count = 26388;
	#10 counter$count = 26389;
	#10 counter$count = 26390;
	#10 counter$count = 26391;
	#10 counter$count = 26392;
	#10 counter$count = 26393;
	#10 counter$count = 26394;
	#10 counter$count = 26395;
	#10 counter$count = 26396;
	#10 counter$count = 26397;
	#10 counter$count = 26398;
	#10 counter$count = 26399;
	#10 counter$count = 26400;
	#10 counter$count = 26401;
	#10 counter$count = 26402;
	#10 counter$count = 26403;
	#10 counter$count = 26404;
	#10 counter$count = 26405;
	#10 counter$count = 26406;
	#10 counter$count = 26407;
	#10 counter$count = 26408;
	#10 counter$count = 26409;
	#10 counter$count = 26410;
	#10 counter$count = 26411;
	#10 counter$count = 26412;
	#10 counter$count = 26413;
	#10 counter$count = 26414;
	#10 counter$count = 26415;
	#10 counter$count = 26416;
	#10 counter$count = 26417;
	#10 counter$count = 26418;
	#10 counter$count = 26419;
	#10 counter$count = 26420;
	#10 counter$count = 26421;
	#10 counter$count = 26422;
	#10 counter$count = 26423;
	#10 counter$count = 26424;
	#10 counter$count = 26425;
	#10 counter$count = 26426;
	#10 counter$count = 26427;
	#10 counter$count = 26428;
	#10 counter$count = 26429;
	#10 counter$count = 26430;
	#10 counter$count = 26431;
	#10 counter$count = 26432;
	#10 counter$count = 26433;
	#10 counter$count = 26434;
	#10 counter$count = 26435;
	#10 counter$count = 26436;
	#10 counter$count = 26437;
	#10 counter$count = 26438;
	#10 counter$count = 26439;
	#10 counter$count = 26440;
	#10 counter$count = 26441;
	#10 counter$count = 26442;
	#10 counter$count = 26443;
	#10 counter$count = 26444;
	#10 counter$count = 26445;
	#10 counter$count = 26446;
	#10 counter$count = 26447;
	#10 counter$count = 26448;
	#10 counter$count = 26449;
	#10 counter$count = 26450;
	#10 counter$count = 26451;
	#10 counter$count = 26452;
	#10 counter$count = 26453;
	#10 counter$count = 26454;
	#10 counter$count = 26455;
	#10 counter$count = 26456;
	#10 counter$count = 26457;
	#10 counter$count = 26458;
	#10 counter$count = 26459;
	#10 counter$count = 26460;
	#10 counter$count = 26461;
	#10 counter$count = 26462;
	#10 counter$count = 26463;
	#10 counter$count = 26464;
	#10 counter$count = 26465;
	#10 counter$count = 26466;
	#10 counter$count = 26467;
	#10 counter$count = 26468;
	#10 counter$count = 26469;
	#10 counter$count = 26470;
	#10 counter$count = 26471;
	#10 counter$count = 26472;
	#10 counter$count = 26473;
	#10 counter$count = 26474;
	#10 counter$count = 26475;
	#10 counter$count = 26476;
	#10 counter$count = 26477;
	#10 counter$count = 26478;
	#10 counter$count = 26479;
	#10 counter$count = 26480;
	#10 counter$count = 26481;
	#10 counter$count = 26482;
	#10 counter$count = 26483;
	#10 counter$count = 26484;
	#10 counter$count = 26485;
	#10 counter$count = 26486;
	#10 counter$count = 26487;
	#10 counter$count = 26488;
	#10 counter$count = 26489;
	#10 counter$count = 26490;
	#10 counter$count = 26491;
	#10 counter$count = 26492;
	#10 counter$count = 26493;
	#10 counter$count = 26494;
	#10 counter$count = 26495;
	#10 counter$count = 26496;
	#10 counter$count = 26497;
	#10 counter$count = 26498;
	#10 counter$count = 26499;
	#10 counter$count = 26500;
	#10 counter$count = 26501;
	#10 counter$count = 26502;
	#10 counter$count = 26503;
	#10 counter$count = 26504;
	#10 counter$count = 26505;
	#10 counter$count = 26506;
	#10 counter$count = 26507;
	#10 counter$count = 26508;
	#10 counter$count = 26509;
	#10 counter$count = 26510;
	#10 counter$count = 26511;
	#10 counter$count = 26512;
	#10 counter$count = 26513;
	#10 counter$count = 26514;
	#10 counter$count = 26515;
	#10 counter$count = 26516;
	#10 counter$count = 26517;
	#10 counter$count = 26518;
	#10 counter$count = 26519;
	#10 counter$count = 26520;
	#10 counter$count = 26521;
	#10 counter$count = 26522;
	#10 counter$count = 26523;
	#10 counter$count = 26524;
	#10 counter$count = 26525;
	#10 counter$count = 26526;
	#10 counter$count = 26527;
	#10 counter$count = 26528;
	#10 counter$count = 26529;
	#10 counter$count = 26530;
	#10 counter$count = 26531;
	#10 counter$count = 26532;
	#10 counter$count = 26533;
	#10 counter$count = 26534;
	#10 counter$count = 26535;
	#10 counter$count = 26536;
	#10 counter$count = 26537;
	#10 counter$count = 26538;
	#10 counter$count = 26539;
	#10 counter$count = 26540;
	#10 counter$count = 26541;
	#10 counter$count = 26542;
	#10 counter$count = 26543;
	#10 counter$count = 26544;
	#10 counter$count = 26545;
	#10 counter$count = 26546;
	#10 counter$count = 26547;
	#10 counter$count = 26548;
	#10 counter$count = 26549;
	#10 counter$count = 26550;
	#10 counter$count = 26551;
	#10 counter$count = 26552;
	#10 counter$count = 26553;
	#10 counter$count = 26554;
	#10 counter$count = 26555;
	#10 counter$count = 26556;
	#10 counter$count = 26557;
	#10 counter$count = 26558;
	#10 counter$count = 26559;
	#10 counter$count = 26560;
	#10 counter$count = 26561;
	#10 counter$count = 26562;
	#10 counter$count = 26563;
	#10 counter$count = 26564;
	#10 counter$count = 26565;
	#10 counter$count = 26566;
	#10 counter$count = 26567;
	#10 counter$count = 26568;
	#10 counter$count = 26569;
	#10 counter$count = 26570;
	#10 counter$count = 26571;
	#10 counter$count = 26572;
	#10 counter$count = 26573;
	#10 counter$count = 26574;
	#10 counter$count = 26575;
	#10 counter$count = 26576;
	#10 counter$count = 26577;
	#10 counter$count = 26578;
	#10 counter$count = 26579;
	#10 counter$count = 26580;
	#10 counter$count = 26581;
	#10 counter$count = 26582;
	#10 counter$count = 26583;
	#10 counter$count = 26584;
	#10 counter$count = 26585;
	#10 counter$count = 26586;
	#10 counter$count = 26587;
	#10 counter$count = 26588;
	#10 counter$count = 26589;
	#10 counter$count = 26590;
	#10 counter$count = 26591;
	#10 counter$count = 26592;
	#10 counter$count = 26593;
	#10 counter$count = 26594;
	#10 counter$count = 26595;
	#10 counter$count = 26596;
	#10 counter$count = 26597;
	#10 counter$count = 26598;
	#10 counter$count = 26599;
	#10 counter$count = 26600;
	#10 counter$count = 26601;
	#10 counter$count = 26602;
	#10 counter$count = 26603;
	#10 counter$count = 26604;
	#10 counter$count = 26605;
	#10 counter$count = 26606;
	#10 counter$count = 26607;
	#10 counter$count = 26608;
	#10 counter$count = 26609;
	#10 counter$count = 26610;
	#10 counter$count = 26611;
	#10 counter$count = 26612;
	#10 counter$count = 26613;
	#10 counter$count = 26614;
	#10 counter$count = 26615;
	#10 counter$count = 26616;
	#10 counter$count = 26617;
	#10 counter$count = 26618;
	#10 counter$count = 26619;
	#10 counter$count = 26620;
	#10 counter$count = 26621;
	#10 counter$count = 26622;
	#10 counter$count = 26623;
	#10 counter$count = 26624;
	#10 counter$count = 26625;
	#10 counter$count = 26626;
	#10 counter$count = 26627;
	#10 counter$count = 26628;
	#10 counter$count = 26629;
	#10 counter$count = 26630;
	#10 counter$count = 26631;
	#10 counter$count = 26632;
	#10 counter$count = 26633;
	#10 counter$count = 26634;
	#10 counter$count = 26635;
	#10 counter$count = 26636;
	#10 counter$count = 26637;
	#10 counter$count = 26638;
	#10 counter$count = 26639;
	#10 counter$count = 26640;
	#10 counter$count = 26641;
	#10 counter$count = 26642;
	#10 counter$count = 26643;
	#10 counter$count = 26644;
	#10 counter$count = 26645;
	#10 counter$count = 26646;
	#10 counter$count = 26647;
	#10 counter$count = 26648;
	#10 counter$count = 26649;
	#10 counter$count = 26650;
	#10 counter$count = 26651;
	#10 counter$count = 26652;
	#10 counter$count = 26653;
	#10 counter$count = 26654;
	#10 counter$count = 26655;
	#10 counter$count = 26656;
	#10 counter$count = 26657;
	#10 counter$count = 26658;
	#10 counter$count = 26659;
	#10 counter$count = 26660;
	#10 counter$count = 26661;
	#10 counter$count = 26662;
	#10 counter$count = 26663;
	#10 counter$count = 26664;
	#10 counter$count = 26665;
	#10 counter$count = 26666;
	#10 counter$count = 26667;
	#10 counter$count = 26668;
	#10 counter$count = 26669;
	#10 counter$count = 26670;
	#10 counter$count = 26671;
	#10 counter$count = 26672;
	#10 counter$count = 26673;
	#10 counter$count = 26674;
	#10 counter$count = 26675;
	#10 counter$count = 26676;
	#10 counter$count = 26677;
	#10 counter$count = 26678;
	#10 counter$count = 26679;
	#10 counter$count = 26680;
	#10 counter$count = 26681;
	#10 counter$count = 26682;
	#10 counter$count = 26683;
	#10 counter$count = 26684;
	#10 counter$count = 26685;
	#10 counter$count = 26686;
	#10 counter$count = 26687;
	#10 counter$count = 26688;
	#10 counter$count = 26689;
	#10 counter$count = 26690;
	#10 counter$count = 26691;
	#10 counter$count = 26692;
	#10 counter$count = 26693;
	#10 counter$count = 26694;
	#10 counter$count = 26695;
	#10 counter$count = 26696;
	#10 counter$count = 26697;
	#10 counter$count = 26698;
	#10 counter$count = 26699;
	#10 counter$count = 26700;
	#10 counter$count = 26701;
	#10 counter$count = 26702;
	#10 counter$count = 26703;
	#10 counter$count = 26704;
	#10 counter$count = 26705;
	#10 counter$count = 26706;
	#10 counter$count = 26707;
	#10 counter$count = 26708;
	#10 counter$count = 26709;
	#10 counter$count = 26710;
	#10 counter$count = 26711;
	#10 counter$count = 26712;
	#10 counter$count = 26713;
	#10 counter$count = 26714;
	#10 counter$count = 26715;
	#10 counter$count = 26716;
	#10 counter$count = 26717;
	#10 counter$count = 26718;
	#10 counter$count = 26719;
	#10 counter$count = 26720;
	#10 counter$count = 26721;
	#10 counter$count = 26722;
	#10 counter$count = 26723;
	#10 counter$count = 26724;
	#10 counter$count = 26725;
	#10 counter$count = 26726;
	#10 counter$count = 26727;
	#10 counter$count = 26728;
	#10 counter$count = 26729;
	#10 counter$count = 26730;
	#10 counter$count = 26731;
	#10 counter$count = 26732;
	#10 counter$count = 26733;
	#10 counter$count = 26734;
	#10 counter$count = 26735;
	#10 counter$count = 26736;
	#10 counter$count = 26737;
	#10 counter$count = 26738;
	#10 counter$count = 26739;
	#10 counter$count = 26740;
	#10 counter$count = 26741;
	#10 counter$count = 26742;
	#10 counter$count = 26743;
	#10 counter$count = 26744;
	#10 counter$count = 26745;
	#10 counter$count = 26746;
	#10 counter$count = 26747;
	#10 counter$count = 26748;
	#10 counter$count = 26749;
	#10 counter$count = 26750;
	#10 counter$count = 26751;
	#10 counter$count = 26752;
	#10 counter$count = 26753;
	#10 counter$count = 26754;
	#10 counter$count = 26755;
	#10 counter$count = 26756;
	#10 counter$count = 26757;
	#10 counter$count = 26758;
	#10 counter$count = 26759;
	#10 counter$count = 26760;
	#10 counter$count = 26761;
	#10 counter$count = 26762;
	#10 counter$count = 26763;
	#10 counter$count = 26764;
	#10 counter$count = 26765;
	#10 counter$count = 26766;
	#10 counter$count = 26767;
	#10 counter$count = 26768;
	#10 counter$count = 26769;
	#10 counter$count = 26770;
	#10 counter$count = 26771;
	#10 counter$count = 26772;
	#10 counter$count = 26773;
	#10 counter$count = 26774;
	#10 counter$count = 26775;
	#10 counter$count = 26776;
	#10 counter$count = 26777;
	#10 counter$count = 26778;
	#10 counter$count = 26779;
	#10 counter$count = 26780;
	#10 counter$count = 26781;
	#10 counter$count = 26782;
	#10 counter$count = 26783;
	#10 counter$count = 26784;
	#10 counter$count = 26785;
	#10 counter$count = 26786;
	#10 counter$count = 26787;
	#10 counter$count = 26788;
	#10 counter$count = 26789;
	#10 counter$count = 26790;
	#10 counter$count = 26791;
	#10 counter$count = 26792;
	#10 counter$count = 26793;
	#10 counter$count = 26794;
	#10 counter$count = 26795;
	#10 counter$count = 26796;
	#10 counter$count = 26797;
	#10 counter$count = 26798;
	#10 counter$count = 26799;
	#10 counter$count = 26800;
	#10 counter$count = 26801;
	#10 counter$count = 26802;
	#10 counter$count = 26803;
	#10 counter$count = 26804;
	#10 counter$count = 26805;
	#10 counter$count = 26806;
	#10 counter$count = 26807;
	#10 counter$count = 26808;
	#10 counter$count = 26809;
	#10 counter$count = 26810;
	#10 counter$count = 26811;
	#10 counter$count = 26812;
	#10 counter$count = 26813;
	#10 counter$count = 26814;
	#10 counter$count = 26815;
	#10 counter$count = 26816;
	#10 counter$count = 26817;
	#10 counter$count = 26818;
	#10 counter$count = 26819;
	#10 counter$count = 26820;
	#10 counter$count = 26821;
	#10 counter$count = 26822;
	#10 counter$count = 26823;
	#10 counter$count = 26824;
	#10 counter$count = 26825;
	#10 counter$count = 26826;
	#10 counter$count = 26827;
	#10 counter$count = 26828;
	#10 counter$count = 26829;
	#10 counter$count = 26830;
	#10 counter$count = 26831;
	#10 counter$count = 26832;
	#10 counter$count = 26833;
	#10 counter$count = 26834;
	#10 counter$count = 26835;
	#10 counter$count = 26836;
	#10 counter$count = 26837;
	#10 counter$count = 26838;
	#10 counter$count = 26839;
	#10 counter$count = 26840;
	#10 counter$count = 26841;
	#10 counter$count = 26842;
	#10 counter$count = 26843;
	#10 counter$count = 26844;
	#10 counter$count = 26845;
	#10 counter$count = 26846;
	#10 counter$count = 26847;
	#10 counter$count = 26848;
	#10 counter$count = 26849;
	#10 counter$count = 26850;
	#10 counter$count = 26851;
	#10 counter$count = 26852;
	#10 counter$count = 26853;
	#10 counter$count = 26854;
	#10 counter$count = 26855;
	#10 counter$count = 26856;
	#10 counter$count = 26857;
	#10 counter$count = 26858;
	#10 counter$count = 26859;
	#10 counter$count = 26860;
	#10 counter$count = 26861;
	#10 counter$count = 26862;
	#10 counter$count = 26863;
	#10 counter$count = 26864;
	#10 counter$count = 26865;
	#10 counter$count = 26866;
	#10 counter$count = 26867;
	#10 counter$count = 26868;
	#10 counter$count = 26869;
	#10 counter$count = 26870;
	#10 counter$count = 26871;
	#10 counter$count = 26872;
	#10 counter$count = 26873;
	#10 counter$count = 26874;
	#10 counter$count = 26875;
	#10 counter$count = 26876;
	#10 counter$count = 26877;
	#10 counter$count = 26878;
	#10 counter$count = 26879;
	#10 counter$count = 26880;
	#10 counter$count = 26881;
	#10 counter$count = 26882;
	#10 counter$count = 26883;
	#10 counter$count = 26884;
	#10 counter$count = 26885;
	#10 counter$count = 26886;
	#10 counter$count = 26887;
	#10 counter$count = 26888;
	#10 counter$count = 26889;
	#10 counter$count = 26890;
	#10 counter$count = 26891;
	#10 counter$count = 26892;
	#10 counter$count = 26893;
	#10 counter$count = 26894;
	#10 counter$count = 26895;
	#10 counter$count = 26896;
	#10 counter$count = 26897;
	#10 counter$count = 26898;
	#10 counter$count = 26899;
	#10 counter$count = 26900;
	#10 counter$count = 26901;
	#10 counter$count = 26902;
	#10 counter$count = 26903;
	#10 counter$count = 26904;
	#10 counter$count = 26905;
	#10 counter$count = 26906;
	#10 counter$count = 26907;
	#10 counter$count = 26908;
	#10 counter$count = 26909;
	#10 counter$count = 26910;
	#10 counter$count = 26911;
	#10 counter$count = 26912;
	#10 counter$count = 26913;
	#10 counter$count = 26914;
	#10 counter$count = 26915;
	#10 counter$count = 26916;
	#10 counter$count = 26917;
	#10 counter$count = 26918;
	#10 counter$count = 26919;
	#10 counter$count = 26920;
	#10 counter$count = 26921;
	#10 counter$count = 26922;
	#10 counter$count = 26923;
	#10 counter$count = 26924;
	#10 counter$count = 26925;
	#10 counter$count = 26926;
	#10 counter$count = 26927;
	#10 counter$count = 26928;
	#10 counter$count = 26929;
	#10 counter$count = 26930;
	#10 counter$count = 26931;
	#10 counter$count = 26932;
	#10 counter$count = 26933;
	#10 counter$count = 26934;
	#10 counter$count = 26935;
	#10 counter$count = 26936;
	#10 counter$count = 26937;
	#10 counter$count = 26938;
	#10 counter$count = 26939;
	#10 counter$count = 26940;
	#10 counter$count = 26941;
	#10 counter$count = 26942;
	#10 counter$count = 26943;
	#10 counter$count = 26944;
	#10 counter$count = 26945;
	#10 counter$count = 26946;
	#10 counter$count = 26947;
	#10 counter$count = 26948;
	#10 counter$count = 26949;
	#10 counter$count = 26950;
	#10 counter$count = 26951;
	#10 counter$count = 26952;
	#10 counter$count = 26953;
	#10 counter$count = 26954;
	#10 counter$count = 26955;
	#10 counter$count = 26956;
	#10 counter$count = 26957;
	#10 counter$count = 26958;
	#10 counter$count = 26959;
	#10 counter$count = 26960;
	#10 counter$count = 26961;
	#10 counter$count = 26962;
	#10 counter$count = 26963;
	#10 counter$count = 26964;
	#10 counter$count = 26965;
	#10 counter$count = 26966;
	#10 counter$count = 26967;
	#10 counter$count = 26968;
	#10 counter$count = 26969;
	#10 counter$count = 26970;
	#10 counter$count = 26971;
	#10 counter$count = 26972;
	#10 counter$count = 26973;
	#10 counter$count = 26974;
	#10 counter$count = 26975;
	#10 counter$count = 26976;
	#10 counter$count = 26977;
	#10 counter$count = 26978;
	#10 counter$count = 26979;
	#10 counter$count = 26980;
	#10 counter$count = 26981;
	#10 counter$count = 26982;
	#10 counter$count = 26983;
	#10 counter$count = 26984;
	#10 counter$count = 26985;
	#10 counter$count = 26986;
	#10 counter$count = 26987;
	#10 counter$count = 26988;
	#10 counter$count = 26989;
	#10 counter$count = 26990;
	#10 counter$count = 26991;
	#10 counter$count = 26992;
	#10 counter$count = 26993;
	#10 counter$count = 26994;
	#10 counter$count = 26995;
	#10 counter$count = 26996;
	#10 counter$count = 26997;
	#10 counter$count = 26998;
	#10 counter$count = 26999;
	#10 counter$count = 27000;
	#10 counter$count = 27001;
	#10 counter$count = 27002;
	#10 counter$count = 27003;
	#10 counter$count = 27004;
	#10 counter$count = 27005;
	#10 counter$count = 27006;
	#10 counter$count = 27007;
	#10 counter$count = 27008;
	#10 counter$count = 27009;
	#10 counter$count = 27010;
	#10 counter$count = 27011;
	#10 counter$count = 27012;
	#10 counter$count = 27013;
	#10 counter$count = 27014;
	#10 counter$count = 27015;
	#10 counter$count = 27016;
	#10 counter$count = 27017;
	#10 counter$count = 27018;
	#10 counter$count = 27019;
	#10 counter$count = 27020;
	#10 counter$count = 27021;
	#10 counter$count = 27022;
	#10 counter$count = 27023;
	#10 counter$count = 27024;
	#10 counter$count = 27025;
	#10 counter$count = 27026;
	#10 counter$count = 27027;
	#10 counter$count = 27028;
	#10 counter$count = 27029;
	#10 counter$count = 27030;
	#10 counter$count = 27031;
	#10 counter$count = 27032;
	#10 counter$count = 27033;
	#10 counter$count = 27034;
	#10 counter$count = 27035;
	#10 counter$count = 27036;
	#10 counter$count = 27037;
	#10 counter$count = 27038;
	#10 counter$count = 27039;
	#10 counter$count = 27040;
	#10 counter$count = 27041;
	#10 counter$count = 27042;
	#10 counter$count = 27043;
	#10 counter$count = 27044;
	#10 counter$count = 27045;
	#10 counter$count = 27046;
	#10 counter$count = 27047;
	#10 counter$count = 27048;
	#10 counter$count = 27049;
	#10 counter$count = 27050;
	#10 counter$count = 27051;
	#10 counter$count = 27052;
	#10 counter$count = 27053;
	#10 counter$count = 27054;
	#10 counter$count = 27055;
	#10 counter$count = 27056;
	#10 counter$count = 27057;
	#10 counter$count = 27058;
	#10 counter$count = 27059;
	#10 counter$count = 27060;
	#10 counter$count = 27061;
	#10 counter$count = 27062;
	#10 counter$count = 27063;
	#10 counter$count = 27064;
	#10 counter$count = 27065;
	#10 counter$count = 27066;
	#10 counter$count = 27067;
	#10 counter$count = 27068;
	#10 counter$count = 27069;
	#10 counter$count = 27070;
	#10 counter$count = 27071;
	#10 counter$count = 27072;
	#10 counter$count = 27073;
	#10 counter$count = 27074;
	#10 counter$count = 27075;
	#10 counter$count = 27076;
	#10 counter$count = 27077;
	#10 counter$count = 27078;
	#10 counter$count = 27079;
	#10 counter$count = 27080;
	#10 counter$count = 27081;
	#10 counter$count = 27082;
	#10 counter$count = 27083;
	#10 counter$count = 27084;
	#10 counter$count = 27085;
	#10 counter$count = 27086;
	#10 counter$count = 27087;
	#10 counter$count = 27088;
	#10 counter$count = 27089;
	#10 counter$count = 27090;
	#10 counter$count = 27091;
	#10 counter$count = 27092;
	#10 counter$count = 27093;
	#10 counter$count = 27094;
	#10 counter$count = 27095;
	#10 counter$count = 27096;
	#10 counter$count = 27097;
	#10 counter$count = 27098;
	#10 counter$count = 27099;
	#10 counter$count = 27100;
	#10 counter$count = 27101;
	#10 counter$count = 27102;
	#10 counter$count = 27103;
	#10 counter$count = 27104;
	#10 counter$count = 27105;
	#10 counter$count = 27106;
	#10 counter$count = 27107;
	#10 counter$count = 27108;
	#10 counter$count = 27109;
	#10 counter$count = 27110;
	#10 counter$count = 27111;
	#10 counter$count = 27112;
	#10 counter$count = 27113;
	#10 counter$count = 27114;
	#10 counter$count = 27115;
	#10 counter$count = 27116;
	#10 counter$count = 27117;
	#10 counter$count = 27118;
	#10 counter$count = 27119;
	#10 counter$count = 27120;
	#10 counter$count = 27121;
	#10 counter$count = 27122;
	#10 counter$count = 27123;
	#10 counter$count = 27124;
	#10 counter$count = 27125;
	#10 counter$count = 27126;
	#10 counter$count = 27127;
	#10 counter$count = 27128;
	#10 counter$count = 27129;
	#10 counter$count = 27130;
	#10 counter$count = 27131;
	#10 counter$count = 27132;
	#10 counter$count = 27133;
	#10 counter$count = 27134;
	#10 counter$count = 27135;
	#10 counter$count = 27136;
	#10 counter$count = 27137;
	#10 counter$count = 27138;
	#10 counter$count = 27139;
	#10 counter$count = 27140;
	#10 counter$count = 27141;
	#10 counter$count = 27142;
	#10 counter$count = 27143;
	#10 counter$count = 27144;
	#10 counter$count = 27145;
	#10 counter$count = 27146;
	#10 counter$count = 27147;
	#10 counter$count = 27148;
	#10 counter$count = 27149;
	#10 counter$count = 27150;
	#10 counter$count = 27151;
	#10 counter$count = 27152;
	#10 counter$count = 27153;
	#10 counter$count = 27154;
	#10 counter$count = 27155;
	#10 counter$count = 27156;
	#10 counter$count = 27157;
	#10 counter$count = 27158;
	#10 counter$count = 27159;
	#10 counter$count = 27160;
	#10 counter$count = 27161;
	#10 counter$count = 27162;
	#10 counter$count = 27163;
	#10 counter$count = 27164;
	#10 counter$count = 27165;
	#10 counter$count = 27166;
	#10 counter$count = 27167;
	#10 counter$count = 27168;
	#10 counter$count = 27169;
	#10 counter$count = 27170;
	#10 counter$count = 27171;
	#10 counter$count = 27172;
	#10 counter$count = 27173;
	#10 counter$count = 27174;
	#10 counter$count = 27175;
	#10 counter$count = 27176;
	#10 counter$count = 27177;
	#10 counter$count = 27178;
	#10 counter$count = 27179;
	#10 counter$count = 27180;
	#10 counter$count = 27181;
	#10 counter$count = 27182;
	#10 counter$count = 27183;
	#10 counter$count = 27184;
	#10 counter$count = 27185;
	#10 counter$count = 27186;
	#10 counter$count = 27187;
	#10 counter$count = 27188;
	#10 counter$count = 27189;
	#10 counter$count = 27190;
	#10 counter$count = 27191;
	#10 counter$count = 27192;
	#10 counter$count = 27193;
	#10 counter$count = 27194;
	#10 counter$count = 27195;
	#10 counter$count = 27196;
	#10 counter$count = 27197;
	#10 counter$count = 27198;
	#10 counter$count = 27199;
	#10 counter$count = 27200;
	#10 counter$count = 27201;
	#10 counter$count = 27202;
	#10 counter$count = 27203;
	#10 counter$count = 27204;
	#10 counter$count = 27205;
	#10 counter$count = 27206;
	#10 counter$count = 27207;
	#10 counter$count = 27208;
	#10 counter$count = 27209;
	#10 counter$count = 27210;
	#10 counter$count = 27211;
	#10 counter$count = 27212;
	#10 counter$count = 27213;
	#10 counter$count = 27214;
	#10 counter$count = 27215;
	#10 counter$count = 27216;
	#10 counter$count = 27217;
	#10 counter$count = 27218;
	#10 counter$count = 27219;
	#10 counter$count = 27220;
	#10 counter$count = 27221;
	#10 counter$count = 27222;
	#10 counter$count = 27223;
	#10 counter$count = 27224;
	#10 counter$count = 27225;
	#10 counter$count = 27226;
	#10 counter$count = 27227;
	#10 counter$count = 27228;
	#10 counter$count = 27229;
	#10 counter$count = 27230;
	#10 counter$count = 27231;
	#10 counter$count = 27232;
	#10 counter$count = 27233;
	#10 counter$count = 27234;
	#10 counter$count = 27235;
	#10 counter$count = 27236;
	#10 counter$count = 27237;
	#10 counter$count = 27238;
	#10 counter$count = 27239;
	#10 counter$count = 27240;
	#10 counter$count = 27241;
	#10 counter$count = 27242;
	#10 counter$count = 27243;
	#10 counter$count = 27244;
	#10 counter$count = 27245;
	#10 counter$count = 27246;
	#10 counter$count = 27247;
	#10 counter$count = 27248;
	#10 counter$count = 27249;
	#10 counter$count = 27250;
	#10 counter$count = 27251;
	#10 counter$count = 27252;
	#10 counter$count = 27253;
	#10 counter$count = 27254;
	#10 counter$count = 27255;
	#10 counter$count = 27256;
	#10 counter$count = 27257;
	#10 counter$count = 27258;
	#10 counter$count = 27259;
	#10 counter$count = 27260;
	#10 counter$count = 27261;
	#10 counter$count = 27262;
	#10 counter$count = 27263;
	#10 counter$count = 27264;
	#10 counter$count = 27265;
	#10 counter$count = 27266;
	#10 counter$count = 27267;
	#10 counter$count = 27268;
	#10 counter$count = 27269;
	#10 counter$count = 27270;
	#10 counter$count = 27271;
	#10 counter$count = 27272;
	#10 counter$count = 27273;
	#10 counter$count = 27274;
	#10 counter$count = 27275;
	#10 counter$count = 27276;
	#10 counter$count = 27277;
	#10 counter$count = 27278;
	#10 counter$count = 27279;
	#10 counter$count = 27280;
	#10 counter$count = 27281;
	#10 counter$count = 27282;
	#10 counter$count = 27283;
	#10 counter$count = 27284;
	#10 counter$count = 27285;
	#10 counter$count = 27286;
	#10 counter$count = 27287;
	#10 counter$count = 27288;
	#10 counter$count = 27289;
	#10 counter$count = 27290;
	#10 counter$count = 27291;
	#10 counter$count = 27292;
	#10 counter$count = 27293;
	#10 counter$count = 27294;
	#10 counter$count = 27295;
	#10 counter$count = 27296;
	#10 counter$count = 27297;
	#10 counter$count = 27298;
	#10 counter$count = 27299;
	#10 counter$count = 27300;
	#10 counter$count = 27301;
	#10 counter$count = 27302;
	#10 counter$count = 27303;
	#10 counter$count = 27304;
	#10 counter$count = 27305;
	#10 counter$count = 27306;
	#10 counter$count = 27307;
	#10 counter$count = 27308;
	#10 counter$count = 27309;
	#10 counter$count = 27310;
	#10 counter$count = 27311;
	#10 counter$count = 27312;
	#10 counter$count = 27313;
	#10 counter$count = 27314;
	#10 counter$count = 27315;
	#10 counter$count = 27316;
	#10 counter$count = 27317;
	#10 counter$count = 27318;
	#10 counter$count = 27319;
	#10 counter$count = 27320;
	#10 counter$count = 27321;
	#10 counter$count = 27322;
	#10 counter$count = 27323;
	#10 counter$count = 27324;
	#10 counter$count = 27325;
	#10 counter$count = 27326;
	#10 counter$count = 27327;
	#10 counter$count = 27328;
	#10 counter$count = 27329;
	#10 counter$count = 27330;
	#10 counter$count = 27331;
	#10 counter$count = 27332;
	#10 counter$count = 27333;
	#10 counter$count = 27334;
	#10 counter$count = 27335;
	#10 counter$count = 27336;
	#10 counter$count = 27337;
	#10 counter$count = 27338;
	#10 counter$count = 27339;
	#10 counter$count = 27340;
	#10 counter$count = 27341;
	#10 counter$count = 27342;
	#10 counter$count = 27343;
	#10 counter$count = 27344;
	#10 counter$count = 27345;
	#10 counter$count = 27346;
	#10 counter$count = 27347;
	#10 counter$count = 27348;
	#10 counter$count = 27349;
	#10 counter$count = 27350;
	#10 counter$count = 27351;
	#10 counter$count = 27352;
	#10 counter$count = 27353;
	#10 counter$count = 27354;
	#10 counter$count = 27355;
	#10 counter$count = 27356;
	#10 counter$count = 27357;
	#10 counter$count = 27358;
	#10 counter$count = 27359;
	#10 counter$count = 27360;
	#10 counter$count = 27361;
	#10 counter$count = 27362;
	#10 counter$count = 27363;
	#10 counter$count = 27364;
	#10 counter$count = 27365;
	#10 counter$count = 27366;
	#10 counter$count = 27367;
	#10 counter$count = 27368;
	#10 counter$count = 27369;
	#10 counter$count = 27370;
	#10 counter$count = 27371;
	#10 counter$count = 27372;
	#10 counter$count = 27373;
	#10 counter$count = 27374;
	#10 counter$count = 27375;
	#10 counter$count = 27376;
	#10 counter$count = 27377;
	#10 counter$count = 27378;
	#10 counter$count = 27379;
	#10 counter$count = 27380;
	#10 counter$count = 27381;
	#10 counter$count = 27382;
	#10 counter$count = 27383;
	#10 counter$count = 27384;
	#10 counter$count = 27385;
	#10 counter$count = 27386;
	#10 counter$count = 27387;
	#10 counter$count = 27388;
	#10 counter$count = 27389;
	#10 counter$count = 27390;
	#10 counter$count = 27391;
	#10 counter$count = 27392;
	#10 counter$count = 27393;
	#10 counter$count = 27394;
	#10 counter$count = 27395;
	#10 counter$count = 27396;
	#10 counter$count = 27397;
	#10 counter$count = 27398;
	#10 counter$count = 27399;
	#10 counter$count = 27400;
	#10 counter$count = 27401;
	#10 counter$count = 27402;
	#10 counter$count = 27403;
	#10 counter$count = 27404;
	#10 counter$count = 27405;
	#10 counter$count = 27406;
	#10 counter$count = 27407;
	#10 counter$count = 27408;
	#10 counter$count = 27409;
	#10 counter$count = 27410;
	#10 counter$count = 27411;
	#10 counter$count = 27412;
	#10 counter$count = 27413;
	#10 counter$count = 27414;
	#10 counter$count = 27415;
	#10 counter$count = 27416;
	#10 counter$count = 27417;
	#10 counter$count = 27418;
	#10 counter$count = 27419;
	#10 counter$count = 27420;
	#10 counter$count = 27421;
	#10 counter$count = 27422;
	#10 counter$count = 27423;
	#10 counter$count = 27424;
	#10 counter$count = 27425;
	#10 counter$count = 27426;
	#10 counter$count = 27427;
	#10 counter$count = 27428;
	#10 counter$count = 27429;
	#10 counter$count = 27430;
	#10 counter$count = 27431;
	#10 counter$count = 27432;
	#10 counter$count = 27433;
	#10 counter$count = 27434;
	#10 counter$count = 27435;
	#10 counter$count = 27436;
	#10 counter$count = 27437;
	#10 counter$count = 27438;
	#10 counter$count = 27439;
	#10 counter$count = 27440;
	#10 counter$count = 27441;
	#10 counter$count = 27442;
	#10 counter$count = 27443;
	#10 counter$count = 27444;
	#10 counter$count = 27445;
	#10 counter$count = 27446;
	#10 counter$count = 27447;
	#10 counter$count = 27448;
	#10 counter$count = 27449;
	#10 counter$count = 27450;
	#10 counter$count = 27451;
	#10 counter$count = 27452;
	#10 counter$count = 27453;
	#10 counter$count = 27454;
	#10 counter$count = 27455;
	#10 counter$count = 27456;
	#10 counter$count = 27457;
	#10 counter$count = 27458;
	#10 counter$count = 27459;
	#10 counter$count = 27460;
	#10 counter$count = 27461;
	#10 counter$count = 27462;
	#10 counter$count = 27463;
	#10 counter$count = 27464;
	#10 counter$count = 27465;
	#10 counter$count = 27466;
	#10 counter$count = 27467;
	#10 counter$count = 27468;
	#10 counter$count = 27469;
	#10 counter$count = 27470;
	#10 counter$count = 27471;
	#10 counter$count = 27472;
	#10 counter$count = 27473;
	#10 counter$count = 27474;
	#10 counter$count = 27475;
	#10 counter$count = 27476;
	#10 counter$count = 27477;
	#10 counter$count = 27478;
	#10 counter$count = 27479;
	#10 counter$count = 27480;
	#10 counter$count = 27481;
	#10 counter$count = 27482;
	#10 counter$count = 27483;
	#10 counter$count = 27484;
	#10 counter$count = 27485;
	#10 counter$count = 27486;
	#10 counter$count = 27487;
	#10 counter$count = 27488;
	#10 counter$count = 27489;
	#10 counter$count = 27490;
	#10 counter$count = 27491;
	#10 counter$count = 27492;
	#10 counter$count = 27493;
	#10 counter$count = 27494;
	#10 counter$count = 27495;
	#10 counter$count = 27496;
	#10 counter$count = 27497;
	#10 counter$count = 27498;
	#10 counter$count = 27499;
	#10 counter$count = 27500;
	#10 counter$count = 27501;
	#10 counter$count = 27502;
	#10 counter$count = 27503;
	#10 counter$count = 27504;
	#10 counter$count = 27505;
	#10 counter$count = 27506;
	#10 counter$count = 27507;
	#10 counter$count = 27508;
	#10 counter$count = 27509;
	#10 counter$count = 27510;
	#10 counter$count = 27511;
	#10 counter$count = 27512;
	#10 counter$count = 27513;
	#10 counter$count = 27514;
	#10 counter$count = 27515;
	#10 counter$count = 27516;
	#10 counter$count = 27517;
	#10 counter$count = 27518;
	#10 counter$count = 27519;
	#10 counter$count = 27520;
	#10 counter$count = 27521;
	#10 counter$count = 27522;
	#10 counter$count = 27523;
	#10 counter$count = 27524;
	#10 counter$count = 27525;
	#10 counter$count = 27526;
	#10 counter$count = 27527;
	#10 counter$count = 27528;
	#10 counter$count = 27529;
	#10 counter$count = 27530;
	#10 counter$count = 27531;
	#10 counter$count = 27532;
	#10 counter$count = 27533;
	#10 counter$count = 27534;
	#10 counter$count = 27535;
	#10 counter$count = 27536;
	#10 counter$count = 27537;
	#10 counter$count = 27538;
	#10 counter$count = 27539;
	#10 counter$count = 27540;
	#10 counter$count = 27541;
	#10 counter$count = 27542;
	#10 counter$count = 27543;
	#10 counter$count = 27544;
	#10 counter$count = 27545;
	#10 counter$count = 27546;
	#10 counter$count = 27547;
	#10 counter$count = 27548;
	#10 counter$count = 27549;
	#10 counter$count = 27550;
	#10 counter$count = 27551;
	#10 counter$count = 27552;
	#10 counter$count = 27553;
	#10 counter$count = 27554;
	#10 counter$count = 27555;
	#10 counter$count = 27556;
	#10 counter$count = 27557;
	#10 counter$count = 27558;
	#10 counter$count = 27559;
	#10 counter$count = 27560;
	#10 counter$count = 27561;
	#10 counter$count = 27562;
	#10 counter$count = 27563;
	#10 counter$count = 27564;
	#10 counter$count = 27565;
	#10 counter$count = 27566;
	#10 counter$count = 27567;
	#10 counter$count = 27568;
	#10 counter$count = 27569;
	#10 counter$count = 27570;
	#10 counter$count = 27571;
	#10 counter$count = 27572;
	#10 counter$count = 27573;
	#10 counter$count = 27574;
	#10 counter$count = 27575;
	#10 counter$count = 27576;
	#10 counter$count = 27577;
	#10 counter$count = 27578;
	#10 counter$count = 27579;
	#10 counter$count = 27580;
	#10 counter$count = 27581;
	#10 counter$count = 27582;
	#10 counter$count = 27583;
	#10 counter$count = 27584;
	#10 counter$count = 27585;
	#10 counter$count = 27586;
	#10 counter$count = 27587;
	#10 counter$count = 27588;
	#10 counter$count = 27589;
	#10 counter$count = 27590;
	#10 counter$count = 27591;
	#10 counter$count = 27592;
	#10 counter$count = 27593;
	#10 counter$count = 27594;
	#10 counter$count = 27595;
	#10 counter$count = 27596;
	#10 counter$count = 27597;
	#10 counter$count = 27598;
	#10 counter$count = 27599;
	#10 counter$count = 27600;
	#10 counter$count = 27601;
	#10 counter$count = 27602;
	#10 counter$count = 27603;
	#10 counter$count = 27604;
	#10 counter$count = 27605;
	#10 counter$count = 27606;
	#10 counter$count = 27607;
	#10 counter$count = 27608;
	#10 counter$count = 27609;
	#10 counter$count = 27610;
	#10 counter$count = 27611;
	#10 counter$count = 27612;
	#10 counter$count = 27613;
	#10 counter$count = 27614;
	#10 counter$count = 27615;
	#10 counter$count = 27616;
	#10 counter$count = 27617;
	#10 counter$count = 27618;
	#10 counter$count = 27619;
	#10 counter$count = 27620;
	#10 counter$count = 27621;
	#10 counter$count = 27622;
	#10 counter$count = 27623;
	#10 counter$count = 27624;
	#10 counter$count = 27625;
	#10 counter$count = 27626;
	#10 counter$count = 27627;
	#10 counter$count = 27628;
	#10 counter$count = 27629;
	#10 counter$count = 27630;
	#10 counter$count = 27631;
	#10 counter$count = 27632;
	#10 counter$count = 27633;
	#10 counter$count = 27634;
	#10 counter$count = 27635;
	#10 counter$count = 27636;
	#10 counter$count = 27637;
	#10 counter$count = 27638;
	#10 counter$count = 27639;
	#10 counter$count = 27640;
	#10 counter$count = 27641;
	#10 counter$count = 27642;
	#10 counter$count = 27643;
	#10 counter$count = 27644;
	#10 counter$count = 27645;
	#10 counter$count = 27646;
	#10 counter$count = 27647;
	#10 counter$count = 27648;
	#10 counter$count = 27649;
	#10 counter$count = 27650;
	#10 counter$count = 27651;
	#10 counter$count = 27652;
	#10 counter$count = 27653;
	#10 counter$count = 27654;
	#10 counter$count = 27655;
	#10 counter$count = 27656;
	#10 counter$count = 27657;
	#10 counter$count = 27658;
	#10 counter$count = 27659;
	#10 counter$count = 27660;
	#10 counter$count = 27661;
	#10 counter$count = 27662;
	#10 counter$count = 27663;
	#10 counter$count = 27664;
	#10 counter$count = 27665;
	#10 counter$count = 27666;
	#10 counter$count = 27667;
	#10 counter$count = 27668;
	#10 counter$count = 27669;
	#10 counter$count = 27670;
	#10 counter$count = 27671;
	#10 counter$count = 27672;
	#10 counter$count = 27673;
	#10 counter$count = 27674;
	#10 counter$count = 27675;
	#10 counter$count = 27676;
	#10 counter$count = 27677;
	#10 counter$count = 27678;
	#10 counter$count = 27679;
	#10 counter$count = 27680;
	#10 counter$count = 27681;
	#10 counter$count = 27682;
	#10 counter$count = 27683;
	#10 counter$count = 27684;
	#10 counter$count = 27685;
	#10 counter$count = 27686;
	#10 counter$count = 27687;
	#10 counter$count = 27688;
	#10 counter$count = 27689;
	#10 counter$count = 27690;
	#10 counter$count = 27691;
	#10 counter$count = 27692;
	#10 counter$count = 27693;
	#10 counter$count = 27694;
	#10 counter$count = 27695;
	#10 counter$count = 27696;
	#10 counter$count = 27697;
	#10 counter$count = 27698;
	#10 counter$count = 27699;
	#10 counter$count = 27700;
	#10 counter$count = 27701;
	#10 counter$count = 27702;
	#10 counter$count = 27703;
	#10 counter$count = 27704;
	#10 counter$count = 27705;
	#10 counter$count = 27706;
	#10 counter$count = 27707;
	#10 counter$count = 27708;
	#10 counter$count = 27709;
	#10 counter$count = 27710;
	#10 counter$count = 27711;
	#10 counter$count = 27712;
	#10 counter$count = 27713;
	#10 counter$count = 27714;
	#10 counter$count = 27715;
	#10 counter$count = 27716;
	#10 counter$count = 27717;
	#10 counter$count = 27718;
	#10 counter$count = 27719;
	#10 counter$count = 27720;
	#10 counter$count = 27721;
	#10 counter$count = 27722;
	#10 counter$count = 27723;
	#10 counter$count = 27724;
	#10 counter$count = 27725;
	#10 counter$count = 27726;
	#10 counter$count = 27727;
	#10 counter$count = 27728;
	#10 counter$count = 27729;
	#10 counter$count = 27730;
	#10 counter$count = 27731;
	#10 counter$count = 27732;
	#10 counter$count = 27733;
	#10 counter$count = 27734;
	#10 counter$count = 27735;
	#10 counter$count = 27736;
	#10 counter$count = 27737;
	#10 counter$count = 27738;
	#10 counter$count = 27739;
	#10 counter$count = 27740;
	#10 counter$count = 27741;
	#10 counter$count = 27742;
	#10 counter$count = 27743;
	#10 counter$count = 27744;
	#10 counter$count = 27745;
	#10 counter$count = 27746;
	#10 counter$count = 27747;
	#10 counter$count = 27748;
	#10 counter$count = 27749;
	#10 counter$count = 27750;
	#10 counter$count = 27751;
	#10 counter$count = 27752;
	#10 counter$count = 27753;
	#10 counter$count = 27754;
	#10 counter$count = 27755;
	#10 counter$count = 27756;
	#10 counter$count = 27757;
	#10 counter$count = 27758;
	#10 counter$count = 27759;
	#10 counter$count = 27760;
	#10 counter$count = 27761;
	#10 counter$count = 27762;
	#10 counter$count = 27763;
	#10 counter$count = 27764;
	#10 counter$count = 27765;
	#10 counter$count = 27766;
	#10 counter$count = 27767;
	#10 counter$count = 27768;
	#10 counter$count = 27769;
	#10 counter$count = 27770;
	#10 counter$count = 27771;
	#10 counter$count = 27772;
	#10 counter$count = 27773;
	#10 counter$count = 27774;
	#10 counter$count = 27775;
	#10 counter$count = 27776;
	#10 counter$count = 27777;
	#10 counter$count = 27778;
	#10 counter$count = 27779;
	#10 counter$count = 27780;
	#10 counter$count = 27781;
	#10 counter$count = 27782;
	#10 counter$count = 27783;
	#10 counter$count = 27784;
	#10 counter$count = 27785;
	#10 counter$count = 27786;
	#10 counter$count = 27787;
	#10 counter$count = 27788;
	#10 counter$count = 27789;
	#10 counter$count = 27790;
	#10 counter$count = 27791;
	#10 counter$count = 27792;
	#10 counter$count = 27793;
	#10 counter$count = 27794;
	#10 counter$count = 27795;
	#10 counter$count = 27796;
	#10 counter$count = 27797;
	#10 counter$count = 27798;
	#10 counter$count = 27799;
	#10 counter$count = 27800;
	#10 counter$count = 27801;
	#10 counter$count = 27802;
	#10 counter$count = 27803;
	#10 counter$count = 27804;
	#10 counter$count = 27805;
	#10 counter$count = 27806;
	#10 counter$count = 27807;
	#10 counter$count = 27808;
	#10 counter$count = 27809;
	#10 counter$count = 27810;
	#10 counter$count = 27811;
	#10 counter$count = 27812;
	#10 counter$count = 27813;
	#10 counter$count = 27814;
	#10 counter$count = 27815;
	#10 counter$count = 27816;
	#10 counter$count = 27817;
	#10 counter$count = 27818;
	#10 counter$count = 27819;
	#10 counter$count = 27820;
	#10 counter$count = 27821;
	#10 counter$count = 27822;
	#10 counter$count = 27823;
	#10 counter$count = 27824;
	#10 counter$count = 27825;
	#10 counter$count = 27826;
	#10 counter$count = 27827;
	#10 counter$count = 27828;
	#10 counter$count = 27829;
	#10 counter$count = 27830;
	#10 counter$count = 27831;
	#10 counter$count = 27832;
	#10 counter$count = 27833;
	#10 counter$count = 27834;
	#10 counter$count = 27835;
	#10 counter$count = 27836;
	#10 counter$count = 27837;
	#10 counter$count = 27838;
	#10 counter$count = 27839;
	#10 counter$count = 27840;
	#10 counter$count = 27841;
	#10 counter$count = 27842;
	#10 counter$count = 27843;
	#10 counter$count = 27844;
	#10 counter$count = 27845;
	#10 counter$count = 27846;
	#10 counter$count = 27847;
	#10 counter$count = 27848;
	#10 counter$count = 27849;
	#10 counter$count = 27850;
	#10 counter$count = 27851;
	#10 counter$count = 27852;
	#10 counter$count = 27853;
	#10 counter$count = 27854;
	#10 counter$count = 27855;
	#10 counter$count = 27856;
	#10 counter$count = 27857;
	#10 counter$count = 27858;
	#10 counter$count = 27859;
	#10 counter$count = 27860;
	#10 counter$count = 27861;
	#10 counter$count = 27862;
	#10 counter$count = 27863;
	#10 counter$count = 27864;
	#10 counter$count = 27865;
	#10 counter$count = 27866;
	#10 counter$count = 27867;
	#10 counter$count = 27868;
	#10 counter$count = 27869;
	#10 counter$count = 27870;
	#10 counter$count = 27871;
	#10 counter$count = 27872;
	#10 counter$count = 27873;
	#10 counter$count = 27874;
	#10 counter$count = 27875;
	#10 counter$count = 27876;
	#10 counter$count = 27877;
	#10 counter$count = 27878;
	#10 counter$count = 27879;
	#10 counter$count = 27880;
	#10 counter$count = 27881;
	#10 counter$count = 27882;
	#10 counter$count = 27883;
	#10 counter$count = 27884;
	#10 counter$count = 27885;
	#10 counter$count = 27886;
	#10 counter$count = 27887;
	#10 counter$count = 27888;
	#10 counter$count = 27889;
	#10 counter$count = 27890;
	#10 counter$count = 27891;
	#10 counter$count = 27892;
	#10 counter$count = 27893;
	#10 counter$count = 27894;
	#10 counter$count = 27895;
	#10 counter$count = 27896;
	#10 counter$count = 27897;
	#10 counter$count = 27898;
	#10 counter$count = 27899;
	#10 counter$count = 27900;
	#10 counter$count = 27901;
	#10 counter$count = 27902;
	#10 counter$count = 27903;
	#10 counter$count = 27904;
	#10 counter$count = 27905;
	#10 counter$count = 27906;
	#10 counter$count = 27907;
	#10 counter$count = 27908;
	#10 counter$count = 27909;
	#10 counter$count = 27910;
	#10 counter$count = 27911;
	#10 counter$count = 27912;
	#10 counter$count = 27913;
	#10 counter$count = 27914;
	#10 counter$count = 27915;
	#10 counter$count = 27916;
	#10 counter$count = 27917;
	#10 counter$count = 27918;
	#10 counter$count = 27919;
	#10 counter$count = 27920;
	#10 counter$count = 27921;
	#10 counter$count = 27922;
	#10 counter$count = 27923;
	#10 counter$count = 27924;
	#10 counter$count = 27925;
	#10 counter$count = 27926;
	#10 counter$count = 27927;
	#10 counter$count = 27928;
	#10 counter$count = 27929;
	#10 counter$count = 27930;
	#10 counter$count = 27931;
	#10 counter$count = 27932;
	#10 counter$count = 27933;
	#10 counter$count = 27934;
	#10 counter$count = 27935;
	#10 counter$count = 27936;
	#10 counter$count = 27937;
	#10 counter$count = 27938;
	#10 counter$count = 27939;
	#10 counter$count = 27940;
	#10 counter$count = 27941;
	#10 counter$count = 27942;
	#10 counter$count = 27943;
	#10 counter$count = 27944;
	#10 counter$count = 27945;
	#10 counter$count = 27946;
	#10 counter$count = 27947;
	#10 counter$count = 27948;
	#10 counter$count = 27949;
	#10 counter$count = 27950;
	#10 counter$count = 27951;
	#10 counter$count = 27952;
	#10 counter$count = 27953;
	#10 counter$count = 27954;
	#10 counter$count = 27955;
	#10 counter$count = 27956;
	#10 counter$count = 27957;
	#10 counter$count = 27958;
	#10 counter$count = 27959;
	#10 counter$count = 27960;
	#10 counter$count = 27961;
	#10 counter$count = 27962;
	#10 counter$count = 27963;
	#10 counter$count = 27964;
	#10 counter$count = 27965;
	#10 counter$count = 27966;
	#10 counter$count = 27967;
	#10 counter$count = 27968;
	#10 counter$count = 27969;
	#10 counter$count = 27970;
	#10 counter$count = 27971;
	#10 counter$count = 27972;
	#10 counter$count = 27973;
	#10 counter$count = 27974;
	#10 counter$count = 27975;
	#10 counter$count = 27976;
	#10 counter$count = 27977;
	#10 counter$count = 27978;
	#10 counter$count = 27979;
	#10 counter$count = 27980;
	#10 counter$count = 27981;
	#10 counter$count = 27982;
	#10 counter$count = 27983;
	#10 counter$count = 27984;
	#10 counter$count = 27985;
	#10 counter$count = 27986;
	#10 counter$count = 27987;
	#10 counter$count = 27988;
	#10 counter$count = 27989;
	#10 counter$count = 27990;
	#10 counter$count = 27991;
	#10 counter$count = 27992;
	#10 counter$count = 27993;
	#10 counter$count = 27994;
	#10 counter$count = 27995;
	#10 counter$count = 27996;
	#10 counter$count = 27997;
	#10 counter$count = 27998;
	#10 counter$count = 27999;
	#10 counter$count = 28000;
	#10 counter$count = 28001;
	#10 counter$count = 28002;
	#10 counter$count = 28003;
	#10 counter$count = 28004;
	#10 counter$count = 28005;
	#10 counter$count = 28006;
	#10 counter$count = 28007;
	#10 counter$count = 28008;
	#10 counter$count = 28009;
	#10 counter$count = 28010;
	#10 counter$count = 28011;
	#10 counter$count = 28012;
	#10 counter$count = 28013;
	#10 counter$count = 28014;
	#10 counter$count = 28015;
	#10 counter$count = 28016;
	#10 counter$count = 28017;
	#10 counter$count = 28018;
	#10 counter$count = 28019;
	#10 counter$count = 28020;
	#10 counter$count = 28021;
	#10 counter$count = 28022;
	#10 counter$count = 28023;
	#10 counter$count = 28024;
	#10 counter$count = 28025;
	#10 counter$count = 28026;
	#10 counter$count = 28027;
	#10 counter$count = 28028;
	#10 counter$count = 28029;
	#10 counter$count = 28030;
	#10 counter$count = 28031;
	#10 counter$count = 28032;
	#10 counter$count = 28033;
	#10 counter$count = 28034;
	#10 counter$count = 28035;
	#10 counter$count = 28036;
	#10 counter$count = 28037;
	#10 counter$count = 28038;
	#10 counter$count = 28039;
	#10 counter$count = 28040;
	#10 counter$count = 28041;
	#10 counter$count = 28042;
	#10 counter$count = 28043;
	#10 counter$count = 28044;
	#10 counter$count = 28045;
	#10 counter$count = 28046;
	#10 counter$count = 28047;
	#10 counter$count = 28048;
	#10 counter$count = 28049;
	#10 counter$count = 28050;
	#10 counter$count = 28051;
	#10 counter$count = 28052;
	#10 counter$count = 28053;
	#10 counter$count = 28054;
	#10 counter$count = 28055;
	#10 counter$count = 28056;
	#10 counter$count = 28057;
	#10 counter$count = 28058;
	#10 counter$count = 28059;
	#10 counter$count = 28060;
	#10 counter$count = 28061;
	#10 counter$count = 28062;
	#10 counter$count = 28063;
	#10 counter$count = 28064;
	#10 counter$count = 28065;
	#10 counter$count = 28066;
	#10 counter$count = 28067;
	#10 counter$count = 28068;
	#10 counter$count = 28069;
	#10 counter$count = 28070;
	#10 counter$count = 28071;
	#10 counter$count = 28072;
	#10 counter$count = 28073;
	#10 counter$count = 28074;
	#10 counter$count = 28075;
	#10 counter$count = 28076;
	#10 counter$count = 28077;
	#10 counter$count = 28078;
	#10 counter$count = 28079;
	#10 counter$count = 28080;
	#10 counter$count = 28081;
	#10 counter$count = 28082;
	#10 counter$count = 28083;
	#10 counter$count = 28084;
	#10 counter$count = 28085;
	#10 counter$count = 28086;
	#10 counter$count = 28087;
	#10 counter$count = 28088;
	#10 counter$count = 28089;
	#10 counter$count = 28090;
	#10 counter$count = 28091;
	#10 counter$count = 28092;
	#10 counter$count = 28093;
	#10 counter$count = 28094;
	#10 counter$count = 28095;
	#10 counter$count = 28096;
	#10 counter$count = 28097;
	#10 counter$count = 28098;
	#10 counter$count = 28099;
	#10 counter$count = 28100;
	#10 counter$count = 28101;
	#10 counter$count = 28102;
	#10 counter$count = 28103;
	#10 counter$count = 28104;
	#10 counter$count = 28105;
	#10 counter$count = 28106;
	#10 counter$count = 28107;
	#10 counter$count = 28108;
	#10 counter$count = 28109;
	#10 counter$count = 28110;
	#10 counter$count = 28111;
	#10 counter$count = 28112;
	#10 counter$count = 28113;
	#10 counter$count = 28114;
	#10 counter$count = 28115;
	#10 counter$count = 28116;
	#10 counter$count = 28117;
	#10 counter$count = 28118;
	#10 counter$count = 28119;
	#10 counter$count = 28120;
	#10 counter$count = 28121;
	#10 counter$count = 28122;
	#10 counter$count = 28123;
	#10 counter$count = 28124;
	#10 counter$count = 28125;
	#10 counter$count = 28126;
	#10 counter$count = 28127;
	#10 counter$count = 28128;
	#10 counter$count = 28129;
	#10 counter$count = 28130;
	#10 counter$count = 28131;
	#10 counter$count = 28132;
	#10 counter$count = 28133;
	#10 counter$count = 28134;
	#10 counter$count = 28135;
	#10 counter$count = 28136;
	#10 counter$count = 28137;
	#10 counter$count = 28138;
	#10 counter$count = 28139;
	#10 counter$count = 28140;
	#10 counter$count = 28141;
	#10 counter$count = 28142;
	#10 counter$count = 28143;
	#10 counter$count = 28144;
	#10 counter$count = 28145;
	#10 counter$count = 28146;
	#10 counter$count = 28147;
	#10 counter$count = 28148;
	#10 counter$count = 28149;
	#10 counter$count = 28150;
	#10 counter$count = 28151;
	#10 counter$count = 28152;
	#10 counter$count = 28153;
	#10 counter$count = 28154;
	#10 counter$count = 28155;
	#10 counter$count = 28156;
	#10 counter$count = 28157;
	#10 counter$count = 28158;
	#10 counter$count = 28159;
	#10 counter$count = 28160;
	#10 counter$count = 28161;
	#10 counter$count = 28162;
	#10 counter$count = 28163;
	#10 counter$count = 28164;
	#10 counter$count = 28165;
	#10 counter$count = 28166;
	#10 counter$count = 28167;
	#10 counter$count = 28168;
	#10 counter$count = 28169;
	#10 counter$count = 28170;
	#10 counter$count = 28171;
	#10 counter$count = 28172;
	#10 counter$count = 28173;
	#10 counter$count = 28174;
	#10 counter$count = 28175;
	#10 counter$count = 28176;
	#10 counter$count = 28177;
	#10 counter$count = 28178;
	#10 counter$count = 28179;
	#10 counter$count = 28180;
	#10 counter$count = 28181;
	#10 counter$count = 28182;
	#10 counter$count = 28183;
	#10 counter$count = 28184;
	#10 counter$count = 28185;
	#10 counter$count = 28186;
	#10 counter$count = 28187;
	#10 counter$count = 28188;
	#10 counter$count = 28189;
	#10 counter$count = 28190;
	#10 counter$count = 28191;
	#10 counter$count = 28192;
	#10 counter$count = 28193;
	#10 counter$count = 28194;
	#10 counter$count = 28195;
	#10 counter$count = 28196;
	#10 counter$count = 28197;
	#10 counter$count = 28198;
	#10 counter$count = 28199;
	#10 counter$count = 28200;
	#10 counter$count = 28201;
	#10 counter$count = 28202;
	#10 counter$count = 28203;
	#10 counter$count = 28204;
	#10 counter$count = 28205;
	#10 counter$count = 28206;
	#10 counter$count = 28207;
	#10 counter$count = 28208;
	#10 counter$count = 28209;
	#10 counter$count = 28210;
	#10 counter$count = 28211;
	#10 counter$count = 28212;
	#10 counter$count = 28213;
	#10 counter$count = 28214;
	#10 counter$count = 28215;
	#10 counter$count = 28216;
	#10 counter$count = 28217;
	#10 counter$count = 28218;
	#10 counter$count = 28219;
	#10 counter$count = 28220;
	#10 counter$count = 28221;
	#10 counter$count = 28222;
	#10 counter$count = 28223;
	#10 counter$count = 28224;
	#10 counter$count = 28225;
	#10 counter$count = 28226;
	#10 counter$count = 28227;
	#10 counter$count = 28228;
	#10 counter$count = 28229;
	#10 counter$count = 28230;
	#10 counter$count = 28231;
	#10 counter$count = 28232;
	#10 counter$count = 28233;
	#10 counter$count = 28234;
	#10 counter$count = 28235;
	#10 counter$count = 28236;
	#10 counter$count = 28237;
	#10 counter$count = 28238;
	#10 counter$count = 28239;
	#10 counter$count = 28240;
	#10 counter$count = 28241;
	#10 counter$count = 28242;
	#10 counter$count = 28243;
	#10 counter$count = 28244;
	#10 counter$count = 28245;
	#10 counter$count = 28246;
	#10 counter$count = 28247;
	#10 counter$count = 28248;
	#10 counter$count = 28249;
	#10 counter$count = 28250;
	#10 counter$count = 28251;
	#10 counter$count = 28252;
	#10 counter$count = 28253;
	#10 counter$count = 28254;
	#10 counter$count = 28255;
	#10 counter$count = 28256;
	#10 counter$count = 28257;
	#10 counter$count = 28258;
	#10 counter$count = 28259;
	#10 counter$count = 28260;
	#10 counter$count = 28261;
	#10 counter$count = 28262;
	#10 counter$count = 28263;
	#10 counter$count = 28264;
	#10 counter$count = 28265;
	#10 counter$count = 28266;
	#10 counter$count = 28267;
	#10 counter$count = 28268;
	#10 counter$count = 28269;
	#10 counter$count = 28270;
	#10 counter$count = 28271;
	#10 counter$count = 28272;
	#10 counter$count = 28273;
	#10 counter$count = 28274;
	#10 counter$count = 28275;
	#10 counter$count = 28276;
	#10 counter$count = 28277;
	#10 counter$count = 28278;
	#10 counter$count = 28279;
	#10 counter$count = 28280;
	#10 counter$count = 28281;
	#10 counter$count = 28282;
	#10 counter$count = 28283;
	#10 counter$count = 28284;
	#10 counter$count = 28285;
	#10 counter$count = 28286;
	#10 counter$count = 28287;
	#10 counter$count = 28288;
	#10 counter$count = 28289;
	#10 counter$count = 28290;
	#10 counter$count = 28291;
	#10 counter$count = 28292;
	#10 counter$count = 28293;
	#10 counter$count = 28294;
	#10 counter$count = 28295;
	#10 counter$count = 28296;
	#10 counter$count = 28297;
	#10 counter$count = 28298;
	#10 counter$count = 28299;
	#10 counter$count = 28300;
	#10 counter$count = 28301;
	#10 counter$count = 28302;
	#10 counter$count = 28303;
	#10 counter$count = 28304;
	#10 counter$count = 28305;
	#10 counter$count = 28306;
	#10 counter$count = 28307;
	#10 counter$count = 28308;
	#10 counter$count = 28309;
	#10 counter$count = 28310;
	#10 counter$count = 28311;
	#10 counter$count = 28312;
	#10 counter$count = 28313;
	#10 counter$count = 28314;
	#10 counter$count = 28315;
	#10 counter$count = 28316;
	#10 counter$count = 28317;
	#10 counter$count = 28318;
	#10 counter$count = 28319;
	#10 counter$count = 28320;
	#10 counter$count = 28321;
	#10 counter$count = 28322;
	#10 counter$count = 28323;
	#10 counter$count = 28324;
	#10 counter$count = 28325;
	#10 counter$count = 28326;
	#10 counter$count = 28327;
	#10 counter$count = 28328;
	#10 counter$count = 28329;
	#10 counter$count = 28330;
	#10 counter$count = 28331;
	#10 counter$count = 28332;
	#10 counter$count = 28333;
	#10 counter$count = 28334;
	#10 counter$count = 28335;
	#10 counter$count = 28336;
	#10 counter$count = 28337;
	#10 counter$count = 28338;
	#10 counter$count = 28339;
	#10 counter$count = 28340;
	#10 counter$count = 28341;
	#10 counter$count = 28342;
	#10 counter$count = 28343;
	#10 counter$count = 28344;
	#10 counter$count = 28345;
	#10 counter$count = 28346;
	#10 counter$count = 28347;
	#10 counter$count = 28348;
	#10 counter$count = 28349;
	#10 counter$count = 28350;
	#10 counter$count = 28351;
	#10 counter$count = 28352;
	#10 counter$count = 28353;
	#10 counter$count = 28354;
	#10 counter$count = 28355;
	#10 counter$count = 28356;
	#10 counter$count = 28357;
	#10 counter$count = 28358;
	#10 counter$count = 28359;
	#10 counter$count = 28360;
	#10 counter$count = 28361;
	#10 counter$count = 28362;
	#10 counter$count = 28363;
	#10 counter$count = 28364;
	#10 counter$count = 28365;
	#10 counter$count = 28366;
	#10 counter$count = 28367;
	#10 counter$count = 28368;
	#10 counter$count = 28369;
	#10 counter$count = 28370;
	#10 counter$count = 28371;
	#10 counter$count = 28372;
	#10 counter$count = 28373;
	#10 counter$count = 28374;
	#10 counter$count = 28375;
	#10 counter$count = 28376;
	#10 counter$count = 28377;
	#10 counter$count = 28378;
	#10 counter$count = 28379;
	#10 counter$count = 28380;
	#10 counter$count = 28381;
	#10 counter$count = 28382;
	#10 counter$count = 28383;
	#10 counter$count = 28384;
	#10 counter$count = 28385;
	#10 counter$count = 28386;
	#10 counter$count = 28387;
	#10 counter$count = 28388;
	#10 counter$count = 28389;
	#10 counter$count = 28390;
	#10 counter$count = 28391;
	#10 counter$count = 28392;
	#10 counter$count = 28393;
	#10 counter$count = 28394;
	#10 counter$count = 28395;
	#10 counter$count = 28396;
	#10 counter$count = 28397;
	#10 counter$count = 28398;
	#10 counter$count = 28399;
	#10 counter$count = 28400;
	#10 counter$count = 28401;
	#10 counter$count = 28402;
	#10 counter$count = 28403;
	#10 counter$count = 28404;
	#10 counter$count = 28405;
	#10 counter$count = 28406;
	#10 counter$count = 28407;
	#10 counter$count = 28408;
	#10 counter$count = 28409;
	#10 counter$count = 28410;
	#10 counter$count = 28411;
	#10 counter$count = 28412;
	#10 counter$count = 28413;
	#10 counter$count = 28414;
	#10 counter$count = 28415;
	#10 counter$count = 28416;
	#10 counter$count = 28417;
	#10 counter$count = 28418;
	#10 counter$count = 28419;
	#10 counter$count = 28420;
	#10 counter$count = 28421;
	#10 counter$count = 28422;
	#10 counter$count = 28423;
	#10 counter$count = 28424;
	#10 counter$count = 28425;
	#10 counter$count = 28426;
	#10 counter$count = 28427;
	#10 counter$count = 28428;
	#10 counter$count = 28429;
	#10 counter$count = 28430;
	#10 counter$count = 28431;
	#10 counter$count = 28432;
	#10 counter$count = 28433;
	#10 counter$count = 28434;
	#10 counter$count = 28435;
	#10 counter$count = 28436;
	#10 counter$count = 28437;
	#10 counter$count = 28438;
	#10 counter$count = 28439;
	#10 counter$count = 28440;
	#10 counter$count = 28441;
	#10 counter$count = 28442;
	#10 counter$count = 28443;
	#10 counter$count = 28444;
	#10 counter$count = 28445;
	#10 counter$count = 28446;
	#10 counter$count = 28447;
	#10 counter$count = 28448;
	#10 counter$count = 28449;
	#10 counter$count = 28450;
	#10 counter$count = 28451;
	#10 counter$count = 28452;
	#10 counter$count = 28453;
	#10 counter$count = 28454;
	#10 counter$count = 28455;
	#10 counter$count = 28456;
	#10 counter$count = 28457;
	#10 counter$count = 28458;
	#10 counter$count = 28459;
	#10 counter$count = 28460;
	#10 counter$count = 28461;
	#10 counter$count = 28462;
	#10 counter$count = 28463;
	#10 counter$count = 28464;
	#10 counter$count = 28465;
	#10 counter$count = 28466;
	#10 counter$count = 28467;
	#10 counter$count = 28468;
	#10 counter$count = 28469;
	#10 counter$count = 28470;
	#10 counter$count = 28471;
	#10 counter$count = 28472;
	#10 counter$count = 28473;
	#10 counter$count = 28474;
	#10 counter$count = 28475;
	#10 counter$count = 28476;
	#10 counter$count = 28477;
	#10 counter$count = 28478;
	#10 counter$count = 28479;
	#10 counter$count = 28480;
	#10 counter$count = 28481;
	#10 counter$count = 28482;
	#10 counter$count = 28483;
	#10 counter$count = 28484;
	#10 counter$count = 28485;
	#10 counter$count = 28486;
	#10 counter$count = 28487;
	#10 counter$count = 28488;
	#10 counter$count = 28489;
	#10 counter$count = 28490;
	#10 counter$count = 28491;
	#10 counter$count = 28492;
	#10 counter$count = 28493;
	#10 counter$count = 28494;
	#10 counter$count = 28495;
	#10 counter$count = 28496;
	#10 counter$count = 28497;
	#10 counter$count = 28498;
	#10 counter$count = 28499;
	#10 counter$count = 28500;
	#10 counter$count = 28501;
	#10 counter$count = 28502;
	#10 counter$count = 28503;
	#10 counter$count = 28504;
	#10 counter$count = 28505;
	#10 counter$count = 28506;
	#10 counter$count = 28507;
	#10 counter$count = 28508;
	#10 counter$count = 28509;
	#10 counter$count = 28510;
	#10 counter$count = 28511;
	#10 counter$count = 28512;
	#10 counter$count = 28513;
	#10 counter$count = 28514;
	#10 counter$count = 28515;
	#10 counter$count = 28516;
	#10 counter$count = 28517;
	#10 counter$count = 28518;
	#10 counter$count = 28519;
	#10 counter$count = 28520;
	#10 counter$count = 28521;
	#10 counter$count = 28522;
	#10 counter$count = 28523;
	#10 counter$count = 28524;
	#10 counter$count = 28525;
	#10 counter$count = 28526;
	#10 counter$count = 28527;
	#10 counter$count = 28528;
	#10 counter$count = 28529;
	#10 counter$count = 28530;
	#10 counter$count = 28531;
	#10 counter$count = 28532;
	#10 counter$count = 28533;
	#10 counter$count = 28534;
	#10 counter$count = 28535;
	#10 counter$count = 28536;
	#10 counter$count = 28537;
	#10 counter$count = 28538;
	#10 counter$count = 28539;
	#10 counter$count = 28540;
	#10 counter$count = 28541;
	#10 counter$count = 28542;
	#10 counter$count = 28543;
	#10 counter$count = 28544;
	#10 counter$count = 28545;
	#10 counter$count = 28546;
	#10 counter$count = 28547;
	#10 counter$count = 28548;
	#10 counter$count = 28549;
	#10 counter$count = 28550;
	#10 counter$count = 28551;
	#10 counter$count = 28552;
	#10 counter$count = 28553;
	#10 counter$count = 28554;
	#10 counter$count = 28555;
	#10 counter$count = 28556;
	#10 counter$count = 28557;
	#10 counter$count = 28558;
	#10 counter$count = 28559;
	#10 counter$count = 28560;
	#10 counter$count = 28561;
	#10 counter$count = 28562;
	#10 counter$count = 28563;
	#10 counter$count = 28564;
	#10 counter$count = 28565;
	#10 counter$count = 28566;
	#10 counter$count = 28567;
	#10 counter$count = 28568;
	#10 counter$count = 28569;
	#10 counter$count = 28570;
	#10 counter$count = 28571;
	#10 counter$count = 28572;
	#10 counter$count = 28573;
	#10 counter$count = 28574;
	#10 counter$count = 28575;
	#10 counter$count = 28576;
	#10 counter$count = 28577;
	#10 counter$count = 28578;
	#10 counter$count = 28579;
	#10 counter$count = 28580;
	#10 counter$count = 28581;
	#10 counter$count = 28582;
	#10 counter$count = 28583;
	#10 counter$count = 28584;
	#10 counter$count = 28585;
	#10 counter$count = 28586;
	#10 counter$count = 28587;
	#10 counter$count = 28588;
	#10 counter$count = 28589;
	#10 counter$count = 28590;
	#10 counter$count = 28591;
	#10 counter$count = 28592;
	#10 counter$count = 28593;
	#10 counter$count = 28594;
	#10 counter$count = 28595;
	#10 counter$count = 28596;
	#10 counter$count = 28597;
	#10 counter$count = 28598;
	#10 counter$count = 28599;
	#10 counter$count = 28600;
	#10 counter$count = 28601;
	#10 counter$count = 28602;
	#10 counter$count = 28603;
	#10 counter$count = 28604;
	#10 counter$count = 28605;
	#10 counter$count = 28606;
	#10 counter$count = 28607;
	#10 counter$count = 28608;
	#10 counter$count = 28609;
	#10 counter$count = 28610;
	#10 counter$count = 28611;
	#10 counter$count = 28612;
	#10 counter$count = 28613;
	#10 counter$count = 28614;
	#10 counter$count = 28615;
	#10 counter$count = 28616;
	#10 counter$count = 28617;
	#10 counter$count = 28618;
	#10 counter$count = 28619;
	#10 counter$count = 28620;
	#10 counter$count = 28621;
	#10 counter$count = 28622;
	#10 counter$count = 28623;
	#10 counter$count = 28624;
	#10 counter$count = 28625;
	#10 counter$count = 28626;
	#10 counter$count = 28627;
	#10 counter$count = 28628;
	#10 counter$count = 28629;
	#10 counter$count = 28630;
	#10 counter$count = 28631;
	#10 counter$count = 28632;
	#10 counter$count = 28633;
	#10 counter$count = 28634;
	#10 counter$count = 28635;
	#10 counter$count = 28636;
	#10 counter$count = 28637;
	#10 counter$count = 28638;
	#10 counter$count = 28639;
	#10 counter$count = 28640;
	#10 counter$count = 28641;
	#10 counter$count = 28642;
	#10 counter$count = 28643;
	#10 counter$count = 28644;
	#10 counter$count = 28645;
	#10 counter$count = 28646;
	#10 counter$count = 28647;
	#10 counter$count = 28648;
	#10 counter$count = 28649;
	#10 counter$count = 28650;
	#10 counter$count = 28651;
	#10 counter$count = 28652;
	#10 counter$count = 28653;
	#10 counter$count = 28654;
	#10 counter$count = 28655;
	#10 counter$count = 28656;
	#10 counter$count = 28657;
	#10 counter$count = 28658;
	#10 counter$count = 28659;
	#10 counter$count = 28660;
	#10 counter$count = 28661;
	#10 counter$count = 28662;
	#10 counter$count = 28663;
	#10 counter$count = 28664;
	#10 counter$count = 28665;
	#10 counter$count = 28666;
	#10 counter$count = 28667;
	#10 counter$count = 28668;
	#10 counter$count = 28669;
	#10 counter$count = 28670;
	#10 counter$count = 28671;
	#10 counter$count = 28672;
	#10 counter$count = 28673;
	#10 counter$count = 28674;
	#10 counter$count = 28675;
	#10 counter$count = 28676;
	#10 counter$count = 28677;
	#10 counter$count = 28678;
	#10 counter$count = 28679;
	#10 counter$count = 28680;
	#10 counter$count = 28681;
	#10 counter$count = 28682;
	#10 counter$count = 28683;
	#10 counter$count = 28684;
	#10 counter$count = 28685;
	#10 counter$count = 28686;
	#10 counter$count = 28687;
	#10 counter$count = 28688;
	#10 counter$count = 28689;
	#10 counter$count = 28690;
	#10 counter$count = 28691;
	#10 counter$count = 28692;
	#10 counter$count = 28693;
	#10 counter$count = 28694;
	#10 counter$count = 28695;
	#10 counter$count = 28696;
	#10 counter$count = 28697;
	#10 counter$count = 28698;
	#10 counter$count = 28699;
	#10 counter$count = 28700;
	#10 counter$count = 28701;
	#10 counter$count = 28702;
	#10 counter$count = 28703;
	#10 counter$count = 28704;
	#10 counter$count = 28705;
	#10 counter$count = 28706;
	#10 counter$count = 28707;
	#10 counter$count = 28708;
	#10 counter$count = 28709;
	#10 counter$count = 28710;
	#10 counter$count = 28711;
	#10 counter$count = 28712;
	#10 counter$count = 28713;
	#10 counter$count = 28714;
	#10 counter$count = 28715;
	#10 counter$count = 28716;
	#10 counter$count = 28717;
	#10 counter$count = 28718;
	#10 counter$count = 28719;
	#10 counter$count = 28720;
	#10 counter$count = 28721;
	#10 counter$count = 28722;
	#10 counter$count = 28723;
	#10 counter$count = 28724;
	#10 counter$count = 28725;
	#10 counter$count = 28726;
	#10 counter$count = 28727;
	#10 counter$count = 28728;
	#10 counter$count = 28729;
	#10 counter$count = 28730;
	#10 counter$count = 28731;
	#10 counter$count = 28732;
	#10 counter$count = 28733;
	#10 counter$count = 28734;
	#10 counter$count = 28735;
	#10 counter$count = 28736;
	#10 counter$count = 28737;
	#10 counter$count = 28738;
	#10 counter$count = 28739;
	#10 counter$count = 28740;
	#10 counter$count = 28741;
	#10 counter$count = 28742;
	#10 counter$count = 28743;
	#10 counter$count = 28744;
	#10 counter$count = 28745;
	#10 counter$count = 28746;
	#10 counter$count = 28747;
	#10 counter$count = 28748;
	#10 counter$count = 28749;
	#10 counter$count = 28750;
	#10 counter$count = 28751;
	#10 counter$count = 28752;
	#10 counter$count = 28753;
	#10 counter$count = 28754;
	#10 counter$count = 28755;
	#10 counter$count = 28756;
	#10 counter$count = 28757;
	#10 counter$count = 28758;
	#10 counter$count = 28759;
	#10 counter$count = 28760;
	#10 counter$count = 28761;
	#10 counter$count = 28762;
	#10 counter$count = 28763;
	#10 counter$count = 28764;
	#10 counter$count = 28765;
	#10 counter$count = 28766;
	#10 counter$count = 28767;
	#10 counter$count = 28768;
	#10 counter$count = 28769;
	#10 counter$count = 28770;
	#10 counter$count = 28771;
	#10 counter$count = 28772;
	#10 counter$count = 28773;
	#10 counter$count = 28774;
	#10 counter$count = 28775;
	#10 counter$count = 28776;
	#10 counter$count = 28777;
	#10 counter$count = 28778;
	#10 counter$count = 28779;
	#10 counter$count = 28780;
	#10 counter$count = 28781;
	#10 counter$count = 28782;
	#10 counter$count = 28783;
	#10 counter$count = 28784;
	#10 counter$count = 28785;
	#10 counter$count = 28786;
	#10 counter$count = 28787;
	#10 counter$count = 28788;
	#10 counter$count = 28789;
	#10 counter$count = 28790;
	#10 counter$count = 28791;
	#10 counter$count = 28792;
	#10 counter$count = 28793;
	#10 counter$count = 28794;
	#10 counter$count = 28795;
	#10 counter$count = 28796;
	#10 counter$count = 28797;
	#10 counter$count = 28798;
	#10 counter$count = 28799;
	#10 counter$count = 28800;
	#10 counter$count = 28801;
	#10 counter$count = 28802;
	#10 counter$count = 28803;
	#10 counter$count = 28804;
	#10 counter$count = 28805;
	#10 counter$count = 28806;
	#10 counter$count = 28807;
	#10 counter$count = 28808;
	#10 counter$count = 28809;
	#10 counter$count = 28810;
	#10 counter$count = 28811;
	#10 counter$count = 28812;
	#10 counter$count = 28813;
	#10 counter$count = 28814;
	#10 counter$count = 28815;
	#10 counter$count = 28816;
	#10 counter$count = 28817;
	#10 counter$count = 28818;
	#10 counter$count = 28819;
	#10 counter$count = 28820;
	#10 counter$count = 28821;
	#10 counter$count = 28822;
	#10 counter$count = 28823;
	#10 counter$count = 28824;
	#10 counter$count = 28825;
	#10 counter$count = 28826;
	#10 counter$count = 28827;
	#10 counter$count = 28828;
	#10 counter$count = 28829;
	#10 counter$count = 28830;
	#10 counter$count = 28831;
	#10 counter$count = 28832;
	#10 counter$count = 28833;
	#10 counter$count = 28834;
	#10 counter$count = 28835;
	#10 counter$count = 28836;
	#10 counter$count = 28837;
	#10 counter$count = 28838;
	#10 counter$count = 28839;
	#10 counter$count = 28840;
	#10 counter$count = 28841;
	#10 counter$count = 28842;
	#10 counter$count = 28843;
	#10 counter$count = 28844;
	#10 counter$count = 28845;
	#10 counter$count = 28846;
	#10 counter$count = 28847;
	#10 counter$count = 28848;
	#10 counter$count = 28849;
	#10 counter$count = 28850;
	#10 counter$count = 28851;
	#10 counter$count = 28852;
	#10 counter$count = 28853;
	#10 counter$count = 28854;
	#10 counter$count = 28855;
	#10 counter$count = 28856;
	#10 counter$count = 28857;
	#10 counter$count = 28858;
	#10 counter$count = 28859;
	#10 counter$count = 28860;
	#10 counter$count = 28861;
	#10 counter$count = 28862;
	#10 counter$count = 28863;
	#10 counter$count = 28864;
	#10 counter$count = 28865;
	#10 counter$count = 28866;
	#10 counter$count = 28867;
	#10 counter$count = 28868;
	#10 counter$count = 28869;
	#10 counter$count = 28870;
	#10 counter$count = 28871;
	#10 counter$count = 28872;
	#10 counter$count = 28873;
	#10 counter$count = 28874;
	#10 counter$count = 28875;
	#10 counter$count = 28876;
	#10 counter$count = 28877;
	#10 counter$count = 28878;
	#10 counter$count = 28879;
	#10 counter$count = 28880;
	#10 counter$count = 28881;
	#10 counter$count = 28882;
	#10 counter$count = 28883;
	#10 counter$count = 28884;
	#10 counter$count = 28885;
	#10 counter$count = 28886;
	#10 counter$count = 28887;
	#10 counter$count = 28888;
	#10 counter$count = 28889;
	#10 counter$count = 28890;
	#10 counter$count = 28891;
	#10 counter$count = 28892;
	#10 counter$count = 28893;
	#10 counter$count = 28894;
	#10 counter$count = 28895;
	#10 counter$count = 28896;
	#10 counter$count = 28897;
	#10 counter$count = 28898;
	#10 counter$count = 28899;
	#10 counter$count = 28900;
	#10 counter$count = 28901;
	#10 counter$count = 28902;
	#10 counter$count = 28903;
	#10 counter$count = 28904;
	#10 counter$count = 28905;
	#10 counter$count = 28906;
	#10 counter$count = 28907;
	#10 counter$count = 28908;
	#10 counter$count = 28909;
	#10 counter$count = 28910;
	#10 counter$count = 28911;
	#10 counter$count = 28912;
	#10 counter$count = 28913;
	#10 counter$count = 28914;
	#10 counter$count = 28915;
	#10 counter$count = 28916;
	#10 counter$count = 28917;
	#10 counter$count = 28918;
	#10 counter$count = 28919;
	#10 counter$count = 28920;
	#10 counter$count = 28921;
	#10 counter$count = 28922;
	#10 counter$count = 28923;
	#10 counter$count = 28924;
	#10 counter$count = 28925;
	#10 counter$count = 28926;
	#10 counter$count = 28927;
	#10 counter$count = 28928;
	#10 counter$count = 28929;
	#10 counter$count = 28930;
	#10 counter$count = 28931;
	#10 counter$count = 28932;
	#10 counter$count = 28933;
	#10 counter$count = 28934;
	#10 counter$count = 28935;
	#10 counter$count = 28936;
	#10 counter$count = 28937;
	#10 counter$count = 28938;
	#10 counter$count = 28939;
	#10 counter$count = 28940;
	#10 counter$count = 28941;
	#10 counter$count = 28942;
	#10 counter$count = 28943;
	#10 counter$count = 28944;
	#10 counter$count = 28945;
	#10 counter$count = 28946;
	#10 counter$count = 28947;
	#10 counter$count = 28948;
	#10 counter$count = 28949;
	#10 counter$count = 28950;
	#10 counter$count = 28951;
	#10 counter$count = 28952;
	#10 counter$count = 28953;
	#10 counter$count = 28954;
	#10 counter$count = 28955;
	#10 counter$count = 28956;
	#10 counter$count = 28957;
	#10 counter$count = 28958;
	#10 counter$count = 28959;
	#10 counter$count = 28960;
	#10 counter$count = 28961;
	#10 counter$count = 28962;
	#10 counter$count = 28963;
	#10 counter$count = 28964;
	#10 counter$count = 28965;
	#10 counter$count = 28966;
	#10 counter$count = 28967;
	#10 counter$count = 28968;
	#10 counter$count = 28969;
	#10 counter$count = 28970;
	#10 counter$count = 28971;
	#10 counter$count = 28972;
	#10 counter$count = 28973;
	#10 counter$count = 28974;
	#10 counter$count = 28975;
	#10 counter$count = 28976;
	#10 counter$count = 28977;
	#10 counter$count = 28978;
	#10 counter$count = 28979;
	#10 counter$count = 28980;
	#10 counter$count = 28981;
	#10 counter$count = 28982;
	#10 counter$count = 28983;
	#10 counter$count = 28984;
	#10 counter$count = 28985;
	#10 counter$count = 28986;
	#10 counter$count = 28987;
	#10 counter$count = 28988;
	#10 counter$count = 28989;
	#10 counter$count = 28990;
	#10 counter$count = 28991;
	#10 counter$count = 28992;
	#10 counter$count = 28993;
	#10 counter$count = 28994;
	#10 counter$count = 28995;
	#10 counter$count = 28996;
	#10 counter$count = 28997;
	#10 counter$count = 28998;
	#10 counter$count = 28999;
	#10 counter$count = 29000;
	#10 counter$count = 29001;
	#10 counter$count = 29002;
	#10 counter$count = 29003;
	#10 counter$count = 29004;
	#10 counter$count = 29005;
	#10 counter$count = 29006;
	#10 counter$count = 29007;
	#10 counter$count = 29008;
	#10 counter$count = 29009;
	#10 counter$count = 29010;
	#10 counter$count = 29011;
	#10 counter$count = 29012;
	#10 counter$count = 29013;
	#10 counter$count = 29014;
	#10 counter$count = 29015;
	#10 counter$count = 29016;
	#10 counter$count = 29017;
	#10 counter$count = 29018;
	#10 counter$count = 29019;
	#10 counter$count = 29020;
	#10 counter$count = 29021;
	#10 counter$count = 29022;
	#10 counter$count = 29023;
	#10 counter$count = 29024;
	#10 counter$count = 29025;
	#10 counter$count = 29026;
	#10 counter$count = 29027;
	#10 counter$count = 29028;
	#10 counter$count = 29029;
	#10 counter$count = 29030;
	#10 counter$count = 29031;
	#10 counter$count = 29032;
	#10 counter$count = 29033;
	#10 counter$count = 29034;
	#10 counter$count = 29035;
	#10 counter$count = 29036;
	#10 counter$count = 29037;
	#10 counter$count = 29038;
	#10 counter$count = 29039;
	#10 counter$count = 29040;
	#10 counter$count = 29041;
	#10 counter$count = 29042;
	#10 counter$count = 29043;
	#10 counter$count = 29044;
	#10 counter$count = 29045;
	#10 counter$count = 29046;
	#10 counter$count = 29047;
	#10 counter$count = 29048;
	#10 counter$count = 29049;
	#10 counter$count = 29050;
	#10 counter$count = 29051;
	#10 counter$count = 29052;
	#10 counter$count = 29053;
	#10 counter$count = 29054;
	#10 counter$count = 29055;
	#10 counter$count = 29056;
	#10 counter$count = 29057;
	#10 counter$count = 29058;
	#10 counter$count = 29059;
	#10 counter$count = 29060;
	#10 counter$count = 29061;
	#10 counter$count = 29062;
	#10 counter$count = 29063;
	#10 counter$count = 29064;
	#10 counter$count = 29065;
	#10 counter$count = 29066;
	#10 counter$count = 29067;
	#10 counter$count = 29068;
	#10 counter$count = 29069;
	#10 counter$count = 29070;
	#10 counter$count = 29071;
	#10 counter$count = 29072;
	#10 counter$count = 29073;
	#10 counter$count = 29074;
	#10 counter$count = 29075;
	#10 counter$count = 29076;
	#10 counter$count = 29077;
	#10 counter$count = 29078;
	#10 counter$count = 29079;
	#10 counter$count = 29080;
	#10 counter$count = 29081;
	#10 counter$count = 29082;
	#10 counter$count = 29083;
	#10 counter$count = 29084;
	#10 counter$count = 29085;
	#10 counter$count = 29086;
	#10 counter$count = 29087;
	#10 counter$count = 29088;
	#10 counter$count = 29089;
	#10 counter$count = 29090;
	#10 counter$count = 29091;
	#10 counter$count = 29092;
	#10 counter$count = 29093;
	#10 counter$count = 29094;
	#10 counter$count = 29095;
	#10 counter$count = 29096;
	#10 counter$count = 29097;
	#10 counter$count = 29098;
	#10 counter$count = 29099;
	#10 counter$count = 29100;
	#10 counter$count = 29101;
	#10 counter$count = 29102;
	#10 counter$count = 29103;
	#10 counter$count = 29104;
	#10 counter$count = 29105;
	#10 counter$count = 29106;
	#10 counter$count = 29107;
	#10 counter$count = 29108;
	#10 counter$count = 29109;
	#10 counter$count = 29110;
	#10 counter$count = 29111;
	#10 counter$count = 29112;
	#10 counter$count = 29113;
	#10 counter$count = 29114;
	#10 counter$count = 29115;
	#10 counter$count = 29116;
	#10 counter$count = 29117;
	#10 counter$count = 29118;
	#10 counter$count = 29119;
	#10 counter$count = 29120;
	#10 counter$count = 29121;
	#10 counter$count = 29122;
	#10 counter$count = 29123;
	#10 counter$count = 29124;
	#10 counter$count = 29125;
	#10 counter$count = 29126;
	#10 counter$count = 29127;
	#10 counter$count = 29128;
	#10 counter$count = 29129;
	#10 counter$count = 29130;
	#10 counter$count = 29131;
	#10 counter$count = 29132;
	#10 counter$count = 29133;
	#10 counter$count = 29134;
	#10 counter$count = 29135;
	#10 counter$count = 29136;
	#10 counter$count = 29137;
	#10 counter$count = 29138;
	#10 counter$count = 29139;
	#10 counter$count = 29140;
	#10 counter$count = 29141;
	#10 counter$count = 29142;
	#10 counter$count = 29143;
	#10 counter$count = 29144;
	#10 counter$count = 29145;
	#10 counter$count = 29146;
	#10 counter$count = 29147;
	#10 counter$count = 29148;
	#10 counter$count = 29149;
	#10 counter$count = 29150;
	#10 counter$count = 29151;
	#10 counter$count = 29152;
	#10 counter$count = 29153;
	#10 counter$count = 29154;
	#10 counter$count = 29155;
	#10 counter$count = 29156;
	#10 counter$count = 29157;
	#10 counter$count = 29158;
	#10 counter$count = 29159;
	#10 counter$count = 29160;
	#10 counter$count = 29161;
	#10 counter$count = 29162;
	#10 counter$count = 29163;
	#10 counter$count = 29164;
	#10 counter$count = 29165;
	#10 counter$count = 29166;
	#10 counter$count = 29167;
	#10 counter$count = 29168;
	#10 counter$count = 29169;
	#10 counter$count = 29170;
	#10 counter$count = 29171;
	#10 counter$count = 29172;
	#10 counter$count = 29173;
	#10 counter$count = 29174;
	#10 counter$count = 29175;
	#10 counter$count = 29176;
	#10 counter$count = 29177;
	#10 counter$count = 29178;
	#10 counter$count = 29179;
	#10 counter$count = 29180;
	#10 counter$count = 29181;
	#10 counter$count = 29182;
	#10 counter$count = 29183;
	#10 counter$count = 29184;
	#10 counter$count = 29185;
	#10 counter$count = 29186;
	#10 counter$count = 29187;
	#10 counter$count = 29188;
	#10 counter$count = 29189;
	#10 counter$count = 29190;
	#10 counter$count = 29191;
	#10 counter$count = 29192;
	#10 counter$count = 29193;
	#10 counter$count = 29194;
	#10 counter$count = 29195;
	#10 counter$count = 29196;
	#10 counter$count = 29197;
	#10 counter$count = 29198;
	#10 counter$count = 29199;
	#10 counter$count = 29200;
	#10 counter$count = 29201;
	#10 counter$count = 29202;
	#10 counter$count = 29203;
	#10 counter$count = 29204;
	#10 counter$count = 29205;
	#10 counter$count = 29206;
	#10 counter$count = 29207;
	#10 counter$count = 29208;
	#10 counter$count = 29209;
	#10 counter$count = 29210;
	#10 counter$count = 29211;
	#10 counter$count = 29212;
	#10 counter$count = 29213;
	#10 counter$count = 29214;
	#10 counter$count = 29215;
	#10 counter$count = 29216;
	#10 counter$count = 29217;
	#10 counter$count = 29218;
	#10 counter$count = 29219;
	#10 counter$count = 29220;
	#10 counter$count = 29221;
	#10 counter$count = 29222;
	#10 counter$count = 29223;
	#10 counter$count = 29224;
	#10 counter$count = 29225;
	#10 counter$count = 29226;
	#10 counter$count = 29227;
	#10 counter$count = 29228;
	#10 counter$count = 29229;
	#10 counter$count = 29230;
	#10 counter$count = 29231;
	#10 counter$count = 29232;
	#10 counter$count = 29233;
	#10 counter$count = 29234;
	#10 counter$count = 29235;
	#10 counter$count = 29236;
	#10 counter$count = 29237;
	#10 counter$count = 29238;
	#10 counter$count = 29239;
	#10 counter$count = 29240;
	#10 counter$count = 29241;
	#10 counter$count = 29242;
	#10 counter$count = 29243;
	#10 counter$count = 29244;
	#10 counter$count = 29245;
	#10 counter$count = 29246;
	#10 counter$count = 29247;
	#10 counter$count = 29248;
	#10 counter$count = 29249;
	#10 counter$count = 29250;
	#10 counter$count = 29251;
	#10 counter$count = 29252;
	#10 counter$count = 29253;
	#10 counter$count = 29254;
	#10 counter$count = 29255;
	#10 counter$count = 29256;
	#10 counter$count = 29257;
	#10 counter$count = 29258;
	#10 counter$count = 29259;
	#10 counter$count = 29260;
	#10 counter$count = 29261;
	#10 counter$count = 29262;
	#10 counter$count = 29263;
	#10 counter$count = 29264;
	#10 counter$count = 29265;
	#10 counter$count = 29266;
	#10 counter$count = 29267;
	#10 counter$count = 29268;
	#10 counter$count = 29269;
	#10 counter$count = 29270;
	#10 counter$count = 29271;
	#10 counter$count = 29272;
	#10 counter$count = 29273;
	#10 counter$count = 29274;
	#10 counter$count = 29275;
	#10 counter$count = 29276;
	#10 counter$count = 29277;
	#10 counter$count = 29278;
	#10 counter$count = 29279;
	#10 counter$count = 29280;
	#10 counter$count = 29281;
	#10 counter$count = 29282;
	#10 counter$count = 29283;
	#10 counter$count = 29284;
	#10 counter$count = 29285;
	#10 counter$count = 29286;
	#10 counter$count = 29287;
	#10 counter$count = 29288;
	#10 counter$count = 29289;
	#10 counter$count = 29290;
	#10 counter$count = 29291;
	#10 counter$count = 29292;
	#10 counter$count = 29293;
	#10 counter$count = 29294;
	#10 counter$count = 29295;
	#10 counter$count = 29296;
	#10 counter$count = 29297;
	#10 counter$count = 29298;
	#10 counter$count = 29299;
	#10 counter$count = 29300;
	#10 counter$count = 29301;
	#10 counter$count = 29302;
	#10 counter$count = 29303;
	#10 counter$count = 29304;
	#10 counter$count = 29305;
	#10 counter$count = 29306;
	#10 counter$count = 29307;
	#10 counter$count = 29308;
	#10 counter$count = 29309;
	#10 counter$count = 29310;
	#10 counter$count = 29311;
	#10 counter$count = 29312;
	#10 counter$count = 29313;
	#10 counter$count = 29314;
	#10 counter$count = 29315;
	#10 counter$count = 29316;
	#10 counter$count = 29317;
	#10 counter$count = 29318;
	#10 counter$count = 29319;
	#10 counter$count = 29320;
	#10 counter$count = 29321;
	#10 counter$count = 29322;
	#10 counter$count = 29323;
	#10 counter$count = 29324;
	#10 counter$count = 29325;
	#10 counter$count = 29326;
	#10 counter$count = 29327;
	#10 counter$count = 29328;
	#10 counter$count = 29329;
	#10 counter$count = 29330;
	#10 counter$count = 29331;
	#10 counter$count = 29332;
	#10 counter$count = 29333;
	#10 counter$count = 29334;
	#10 counter$count = 29335;
	#10 counter$count = 29336;
	#10 counter$count = 29337;
	#10 counter$count = 29338;
	#10 counter$count = 29339;
	#10 counter$count = 29340;
	#10 counter$count = 29341;
	#10 counter$count = 29342;
	#10 counter$count = 29343;
	#10 counter$count = 29344;
	#10 counter$count = 29345;
	#10 counter$count = 29346;
	#10 counter$count = 29347;
	#10 counter$count = 29348;
	#10 counter$count = 29349;
	#10 counter$count = 29350;
	#10 counter$count = 29351;
	#10 counter$count = 29352;
	#10 counter$count = 29353;
	#10 counter$count = 29354;
	#10 counter$count = 29355;
	#10 counter$count = 29356;
	#10 counter$count = 29357;
	#10 counter$count = 29358;
	#10 counter$count = 29359;
	#10 counter$count = 29360;
	#10 counter$count = 29361;
	#10 counter$count = 29362;
	#10 counter$count = 29363;
	#10 counter$count = 29364;
	#10 counter$count = 29365;
	#10 counter$count = 29366;
	#10 counter$count = 29367;
	#10 counter$count = 29368;
	#10 counter$count = 29369;
	#10 counter$count = 29370;
	#10 counter$count = 29371;
	#10 counter$count = 29372;
	#10 counter$count = 29373;
	#10 counter$count = 29374;
	#10 counter$count = 29375;
	#10 counter$count = 29376;
	#10 counter$count = 29377;
	#10 counter$count = 29378;
	#10 counter$count = 29379;
	#10 counter$count = 29380;
	#10 counter$count = 29381;
	#10 counter$count = 29382;
	#10 counter$count = 29383;
	#10 counter$count = 29384;
	#10 counter$count = 29385;
	#10 counter$count = 29386;
	#10 counter$count = 29387;
	#10 counter$count = 29388;
	#10 counter$count = 29389;
	#10 counter$count = 29390;
	#10 counter$count = 29391;
	#10 counter$count = 29392;
	#10 counter$count = 29393;
	#10 counter$count = 29394;
	#10 counter$count = 29395;
	#10 counter$count = 29396;
	#10 counter$count = 29397;
	#10 counter$count = 29398;
	#10 counter$count = 29399;
	#10 counter$count = 29400;
	#10 counter$count = 29401;
	#10 counter$count = 29402;
	#10 counter$count = 29403;
	#10 counter$count = 29404;
	#10 counter$count = 29405;
	#10 counter$count = 29406;
	#10 counter$count = 29407;
	#10 counter$count = 29408;
	#10 counter$count = 29409;
	#10 counter$count = 29410;
	#10 counter$count = 29411;
	#10 counter$count = 29412;
	#10 counter$count = 29413;
	#10 counter$count = 29414;
	#10 counter$count = 29415;
	#10 counter$count = 29416;
	#10 counter$count = 29417;
	#10 counter$count = 29418;
	#10 counter$count = 29419;
	#10 counter$count = 29420;
	#10 counter$count = 29421;
	#10 counter$count = 29422;
	#10 counter$count = 29423;
	#10 counter$count = 29424;
	#10 counter$count = 29425;
	#10 counter$count = 29426;
	#10 counter$count = 29427;
	#10 counter$count = 29428;
	#10 counter$count = 29429;
	#10 counter$count = 29430;
	#10 counter$count = 29431;
	#10 counter$count = 29432;
	#10 counter$count = 29433;
	#10 counter$count = 29434;
	#10 counter$count = 29435;
	#10 counter$count = 29436;
	#10 counter$count = 29437;
	#10 counter$count = 29438;
	#10 counter$count = 29439;
	#10 counter$count = 29440;
	#10 counter$count = 29441;
	#10 counter$count = 29442;
	#10 counter$count = 29443;
	#10 counter$count = 29444;
	#10 counter$count = 29445;
	#10 counter$count = 29446;
	#10 counter$count = 29447;
	#10 counter$count = 29448;
	#10 counter$count = 29449;
	#10 counter$count = 29450;
	#10 counter$count = 29451;
	#10 counter$count = 29452;
	#10 counter$count = 29453;
	#10 counter$count = 29454;
	#10 counter$count = 29455;
	#10 counter$count = 29456;
	#10 counter$count = 29457;
	#10 counter$count = 29458;
	#10 counter$count = 29459;
	#10 counter$count = 29460;
	#10 counter$count = 29461;
	#10 counter$count = 29462;
	#10 counter$count = 29463;
	#10 counter$count = 29464;
	#10 counter$count = 29465;
	#10 counter$count = 29466;
	#10 counter$count = 29467;
	#10 counter$count = 29468;
	#10 counter$count = 29469;
	#10 counter$count = 29470;
	#10 counter$count = 29471;
	#10 counter$count = 29472;
	#10 counter$count = 29473;
	#10 counter$count = 29474;
	#10 counter$count = 29475;
	#10 counter$count = 29476;
	#10 counter$count = 29477;
	#10 counter$count = 29478;
	#10 counter$count = 29479;
	#10 counter$count = 29480;
	#10 counter$count = 29481;
	#10 counter$count = 29482;
	#10 counter$count = 29483;
	#10 counter$count = 29484;
	#10 counter$count = 29485;
	#10 counter$count = 29486;
	#10 counter$count = 29487;
	#10 counter$count = 29488;
	#10 counter$count = 29489;
	#10 counter$count = 29490;
	#10 counter$count = 29491;
	#10 counter$count = 29492;
	#10 counter$count = 29493;
	#10 counter$count = 29494;
	#10 counter$count = 29495;
	#10 counter$count = 29496;
	#10 counter$count = 29497;
	#10 counter$count = 29498;
	#10 counter$count = 29499;
	#10 counter$count = 29500;
	#10 counter$count = 29501;
	#10 counter$count = 29502;
	#10 counter$count = 29503;
	#10 counter$count = 29504;
	#10 counter$count = 29505;
	#10 counter$count = 29506;
	#10 counter$count = 29507;
	#10 counter$count = 29508;
	#10 counter$count = 29509;
	#10 counter$count = 29510;
	#10 counter$count = 29511;
	#10 counter$count = 29512;
	#10 counter$count = 29513;
	#10 counter$count = 29514;
	#10 counter$count = 29515;
	#10 counter$count = 29516;
	#10 counter$count = 29517;
	#10 counter$count = 29518;
	#10 counter$count = 29519;
	#10 counter$count = 29520;
	#10 counter$count = 29521;
	#10 counter$count = 29522;
	#10 counter$count = 29523;
	#10 counter$count = 29524;
	#10 counter$count = 29525;
	#10 counter$count = 29526;
	#10 counter$count = 29527;
	#10 counter$count = 29528;
	#10 counter$count = 29529;
	#10 counter$count = 29530;
	#10 counter$count = 29531;
	#10 counter$count = 29532;
	#10 counter$count = 29533;
	#10 counter$count = 29534;
	#10 counter$count = 29535;
	#10 counter$count = 29536;
	#10 counter$count = 29537;
	#10 counter$count = 29538;
	#10 counter$count = 29539;
	#10 counter$count = 29540;
	#10 counter$count = 29541;
	#10 counter$count = 29542;
	#10 counter$count = 29543;
	#10 counter$count = 29544;
	#10 counter$count = 29545;
	#10 counter$count = 29546;
	#10 counter$count = 29547;
	#10 counter$count = 29548;
	#10 counter$count = 29549;
	#10 counter$count = 29550;
	#10 counter$count = 29551;
	#10 counter$count = 29552;
	#10 counter$count = 29553;
	#10 counter$count = 29554;
	#10 counter$count = 29555;
	#10 counter$count = 29556;
	#10 counter$count = 29557;
	#10 counter$count = 29558;
	#10 counter$count = 29559;
	#10 counter$count = 29560;
	#10 counter$count = 29561;
	#10 counter$count = 29562;
	#10 counter$count = 29563;
	#10 counter$count = 29564;
	#10 counter$count = 29565;
	#10 counter$count = 29566;
	#10 counter$count = 29567;
	#10 counter$count = 29568;
	#10 counter$count = 29569;
	#10 counter$count = 29570;
	#10 counter$count = 29571;
	#10 counter$count = 29572;
	#10 counter$count = 29573;
	#10 counter$count = 29574;
	#10 counter$count = 29575;
	#10 counter$count = 29576;
	#10 counter$count = 29577;
	#10 counter$count = 29578;
	#10 counter$count = 29579;
	#10 counter$count = 29580;
	#10 counter$count = 29581;
	#10 counter$count = 29582;
	#10 counter$count = 29583;
	#10 counter$count = 29584;
	#10 counter$count = 29585;
	#10 counter$count = 29586;
	#10 counter$count = 29587;
	#10 counter$count = 29588;
	#10 counter$count = 29589;
	#10 counter$count = 29590;
	#10 counter$count = 29591;
	#10 counter$count = 29592;
	#10 counter$count = 29593;
	#10 counter$count = 29594;
	#10 counter$count = 29595;
	#10 counter$count = 29596;
	#10 counter$count = 29597;
	#10 counter$count = 29598;
	#10 counter$count = 29599;
	#10 counter$count = 29600;
	#10 counter$count = 29601;
	#10 counter$count = 29602;
	#10 counter$count = 29603;
	#10 counter$count = 29604;
	#10 counter$count = 29605;
	#10 counter$count = 29606;
	#10 counter$count = 29607;
	#10 counter$count = 29608;
	#10 counter$count = 29609;
	#10 counter$count = 29610;
	#10 counter$count = 29611;
	#10 counter$count = 29612;
	#10 counter$count = 29613;
	#10 counter$count = 29614;
	#10 counter$count = 29615;
	#10 counter$count = 29616;
	#10 counter$count = 29617;
	#10 counter$count = 29618;
	#10 counter$count = 29619;
	#10 counter$count = 29620;
	#10 counter$count = 29621;
	#10 counter$count = 29622;
	#10 counter$count = 29623;
	#10 counter$count = 29624;
	#10 counter$count = 29625;
	#10 counter$count = 29626;
	#10 counter$count = 29627;
	#10 counter$count = 29628;
	#10 counter$count = 29629;
	#10 counter$count = 29630;
	#10 counter$count = 29631;
	#10 counter$count = 29632;
	#10 counter$count = 29633;
	#10 counter$count = 29634;
	#10 counter$count = 29635;
	#10 counter$count = 29636;
	#10 counter$count = 29637;
	#10 counter$count = 29638;
	#10 counter$count = 29639;
	#10 counter$count = 29640;
	#10 counter$count = 29641;
	#10 counter$count = 29642;
	#10 counter$count = 29643;
	#10 counter$count = 29644;
	#10 counter$count = 29645;
	#10 counter$count = 29646;
	#10 counter$count = 29647;
	#10 counter$count = 29648;
	#10 counter$count = 29649;
	#10 counter$count = 29650;
	#10 counter$count = 29651;
	#10 counter$count = 29652;
	#10 counter$count = 29653;
	#10 counter$count = 29654;
	#10 counter$count = 29655;
	#10 counter$count = 29656;
	#10 counter$count = 29657;
	#10 counter$count = 29658;
	#10 counter$count = 29659;
	#10 counter$count = 29660;
	#10 counter$count = 29661;
	#10 counter$count = 29662;
	#10 counter$count = 29663;
	#10 counter$count = 29664;
	#10 counter$count = 29665;
	#10 counter$count = 29666;
	#10 counter$count = 29667;
	#10 counter$count = 29668;
	#10 counter$count = 29669;
	#10 counter$count = 29670;
	#10 counter$count = 29671;
	#10 counter$count = 29672;
	#10 counter$count = 29673;
	#10 counter$count = 29674;
	#10 counter$count = 29675;
	#10 counter$count = 29676;
	#10 counter$count = 29677;
	#10 counter$count = 29678;
	#10 counter$count = 29679;
	#10 counter$count = 29680;
	#10 counter$count = 29681;
	#10 counter$count = 29682;
	#10 counter$count = 29683;
	#10 counter$count = 29684;
	#10 counter$count = 29685;
	#10 counter$count = 29686;
	#10 counter$count = 29687;
	#10 counter$count = 29688;
	#10 counter$count = 29689;
	#10 counter$count = 29690;
	#10 counter$count = 29691;
	#10 counter$count = 29692;
	#10 counter$count = 29693;
	#10 counter$count = 29694;
	#10 counter$count = 29695;
	#10 counter$count = 29696;
	#10 counter$count = 29697;
	#10 counter$count = 29698;
	#10 counter$count = 29699;
	#10 counter$count = 29700;
	#10 counter$count = 29701;
	#10 counter$count = 29702;
	#10 counter$count = 29703;
	#10 counter$count = 29704;
	#10 counter$count = 29705;
	#10 counter$count = 29706;
	#10 counter$count = 29707;
	#10 counter$count = 29708;
	#10 counter$count = 29709;
	#10 counter$count = 29710;
	#10 counter$count = 29711;
	#10 counter$count = 29712;
	#10 counter$count = 29713;
	#10 counter$count = 29714;
	#10 counter$count = 29715;
	#10 counter$count = 29716;
	#10 counter$count = 29717;
	#10 counter$count = 29718;
	#10 counter$count = 29719;
	#10 counter$count = 29720;
	#10 counter$count = 29721;
	#10 counter$count = 29722;
	#10 counter$count = 29723;
	#10 counter$count = 29724;
	#10 counter$count = 29725;
	#10 counter$count = 29726;
	#10 counter$count = 29727;
	#10 counter$count = 29728;
	#10 counter$count = 29729;
	#10 counter$count = 29730;
	#10 counter$count = 29731;
	#10 counter$count = 29732;
	#10 counter$count = 29733;
	#10 counter$count = 29734;
	#10 counter$count = 29735;
	#10 counter$count = 29736;
	#10 counter$count = 29737;
	#10 counter$count = 29738;
	#10 counter$count = 29739;
	#10 counter$count = 29740;
	#10 counter$count = 29741;
	#10 counter$count = 29742;
	#10 counter$count = 29743;
	#10 counter$count = 29744;
	#10 counter$count = 29745;
	#10 counter$count = 29746;
	#10 counter$count = 29747;
	#10 counter$count = 29748;
	#10 counter$count = 29749;
	#10 counter$count = 29750;
	#10 counter$count = 29751;
	#10 counter$count = 29752;
	#10 counter$count = 29753;
	#10 counter$count = 29754;
	#10 counter$count = 29755;
	#10 counter$count = 29756;
	#10 counter$count = 29757;
	#10 counter$count = 29758;
	#10 counter$count = 29759;
	#10 counter$count = 29760;
	#10 counter$count = 29761;
	#10 counter$count = 29762;
	#10 counter$count = 29763;
	#10 counter$count = 29764;
	#10 counter$count = 29765;
	#10 counter$count = 29766;
	#10 counter$count = 29767;
	#10 counter$count = 29768;
	#10 counter$count = 29769;
	#10 counter$count = 29770;
	#10 counter$count = 29771;
	#10 counter$count = 29772;
	#10 counter$count = 29773;
	#10 counter$count = 29774;
	#10 counter$count = 29775;
	#10 counter$count = 29776;
	#10 counter$count = 29777;
	#10 counter$count = 29778;
	#10 counter$count = 29779;
	#10 counter$count = 29780;
	#10 counter$count = 29781;
	#10 counter$count = 29782;
	#10 counter$count = 29783;
	#10 counter$count = 29784;
	#10 counter$count = 29785;
	#10 counter$count = 29786;
	#10 counter$count = 29787;
	#10 counter$count = 29788;
	#10 counter$count = 29789;
	#10 counter$count = 29790;
	#10 counter$count = 29791;
	#10 counter$count = 29792;
	#10 counter$count = 29793;
	#10 counter$count = 29794;
	#10 counter$count = 29795;
	#10 counter$count = 29796;
	#10 counter$count = 29797;
	#10 counter$count = 29798;
	#10 counter$count = 29799;
	#10 counter$count = 29800;
	#10 counter$count = 29801;
	#10 counter$count = 29802;
	#10 counter$count = 29803;
	#10 counter$count = 29804;
	#10 counter$count = 29805;
	#10 counter$count = 29806;
	#10 counter$count = 29807;
	#10 counter$count = 29808;
	#10 counter$count = 29809;
	#10 counter$count = 29810;
	#10 counter$count = 29811;
	#10 counter$count = 29812;
	#10 counter$count = 29813;
	#10 counter$count = 29814;
	#10 counter$count = 29815;
	#10 counter$count = 29816;
	#10 counter$count = 29817;
	#10 counter$count = 29818;
	#10 counter$count = 29819;
	#10 counter$count = 29820;
	#10 counter$count = 29821;
	#10 counter$count = 29822;
	#10 counter$count = 29823;
	#10 counter$count = 29824;
	#10 counter$count = 29825;
	#10 counter$count = 29826;
	#10 counter$count = 29827;
	#10 counter$count = 29828;
	#10 counter$count = 29829;
	#10 counter$count = 29830;
	#10 counter$count = 29831;
	#10 counter$count = 29832;
	#10 counter$count = 29833;
	#10 counter$count = 29834;
	#10 counter$count = 29835;
	#10 counter$count = 29836;
	#10 counter$count = 29837;
	#10 counter$count = 29838;
	#10 counter$count = 29839;
	#10 counter$count = 29840;
	#10 counter$count = 29841;
	#10 counter$count = 29842;
	#10 counter$count = 29843;
	#10 counter$count = 29844;
	#10 counter$count = 29845;
	#10 counter$count = 29846;
	#10 counter$count = 29847;
	#10 counter$count = 29848;
	#10 counter$count = 29849;
	#10 counter$count = 29850;
	#10 counter$count = 29851;
	#10 counter$count = 29852;
	#10 counter$count = 29853;
	#10 counter$count = 29854;
	#10 counter$count = 29855;
	#10 counter$count = 29856;
	#10 counter$count = 29857;
	#10 counter$count = 29858;
	#10 counter$count = 29859;
	#10 counter$count = 29860;
	#10 counter$count = 29861;
	#10 counter$count = 29862;
	#10 counter$count = 29863;
	#10 counter$count = 29864;
	#10 counter$count = 29865;
	#10 counter$count = 29866;
	#10 counter$count = 29867;
	#10 counter$count = 29868;
	#10 counter$count = 29869;
	#10 counter$count = 29870;
	#10 counter$count = 29871;
	#10 counter$count = 29872;
	#10 counter$count = 29873;
	#10 counter$count = 29874;
	#10 counter$count = 29875;
	#10 counter$count = 29876;
	#10 counter$count = 29877;
	#10 counter$count = 29878;
	#10 counter$count = 29879;
	#10 counter$count = 29880;
	#10 counter$count = 29881;
	#10 counter$count = 29882;
	#10 counter$count = 29883;
	#10 counter$count = 29884;
	#10 counter$count = 29885;
	#10 counter$count = 29886;
	#10 counter$count = 29887;
	#10 counter$count = 29888;
	#10 counter$count = 29889;
	#10 counter$count = 29890;
	#10 counter$count = 29891;
	#10 counter$count = 29892;
	#10 counter$count = 29893;
	#10 counter$count = 29894;
	#10 counter$count = 29895;
	#10 counter$count = 29896;
	#10 counter$count = 29897;
	#10 counter$count = 29898;
	#10 counter$count = 29899;
	#10 counter$count = 29900;
	#10 counter$count = 29901;
	#10 counter$count = 29902;
	#10 counter$count = 29903;
	#10 counter$count = 29904;
	#10 counter$count = 29905;
	#10 counter$count = 29906;
	#10 counter$count = 29907;
	#10 counter$count = 29908;
	#10 counter$count = 29909;
	#10 counter$count = 29910;
	#10 counter$count = 29911;
	#10 counter$count = 29912;
	#10 counter$count = 29913;
	#10 counter$count = 29914;
	#10 counter$count = 29915;
	#10 counter$count = 29916;
	#10 counter$count = 29917;
	#10 counter$count = 29918;
	#10 counter$count = 29919;
	#10 counter$count = 29920;
	#10 counter$count = 29921;
	#10 counter$count = 29922;
	#10 counter$count = 29923;
	#10 counter$count = 29924;
	#10 counter$count = 29925;
	#10 counter$count = 29926;
	#10 counter$count = 29927;
	#10 counter$count = 29928;
	#10 counter$count = 29929;
	#10 counter$count = 29930;
	#10 counter$count = 29931;
	#10 counter$count = 29932;
	#10 counter$count = 29933;
	#10 counter$count = 29934;
	#10 counter$count = 29935;
	#10 counter$count = 29936;
	#10 counter$count = 29937;
	#10 counter$count = 29938;
	#10 counter$count = 29939;
	#10 counter$count = 29940;
	#10 counter$count = 29941;
	#10 counter$count = 29942;
	#10 counter$count = 29943;
	#10 counter$count = 29944;
	#10 counter$count = 29945;
	#10 counter$count = 29946;
	#10 counter$count = 29947;
	#10 counter$count = 29948;
	#10 counter$count = 29949;
	#10 counter$count = 29950;
	#10 counter$count = 29951;
	#10 counter$count = 29952;
	#10 counter$count = 29953;
	#10 counter$count = 29954;
	#10 counter$count = 29955;
	#10 counter$count = 29956;
	#10 counter$count = 29957;
	#10 counter$count = 29958;
	#10 counter$count = 29959;
	#10 counter$count = 29960;
	#10 counter$count = 29961;
	#10 counter$count = 29962;
	#10 counter$count = 29963;
	#10 counter$count = 29964;
	#10 counter$count = 29965;
	#10 counter$count = 29966;
	#10 counter$count = 29967;
	#10 counter$count = 29968;
	#10 counter$count = 29969;
	#10 counter$count = 29970;
	#10 counter$count = 29971;
	#10 counter$count = 29972;
	#10 counter$count = 29973;
	#10 counter$count = 29974;
	#10 counter$count = 29975;
	#10 counter$count = 29976;
	#10 counter$count = 29977;
	#10 counter$count = 29978;
	#10 counter$count = 29979;
	#10 counter$count = 29980;
	#10 counter$count = 29981;
	#10 counter$count = 29982;
	#10 counter$count = 29983;
	#10 counter$count = 29984;
	#10 counter$count = 29985;
	#10 counter$count = 29986;
	#10 counter$count = 29987;
	#10 counter$count = 29988;
	#10 counter$count = 29989;
	#10 counter$count = 29990;
	#10 counter$count = 29991;
	#10 counter$count = 29992;
	#10 counter$count = 29993;
	#10 counter$count = 29994;
	#10 counter$count = 29995;
	#10 counter$count = 29996;
	#10 counter$count = 29997;
	#10 counter$count = 29998;
	#10 counter$count = 29999;
	#10 counter$count = 30000;
	#10 counter$count = 30001;
	#10 counter$count = 30002;
	#10 counter$count = 30003;
	#10 counter$count = 30004;
	#10 counter$count = 30005;
	#10 counter$count = 30006;
	#10 counter$count = 30007;
	#10 counter$count = 30008;
	#10 counter$count = 30009;
	#10 counter$count = 30010;
	#10 counter$count = 30011;
	#10 counter$count = 30012;
	#10 counter$count = 30013;
	#10 counter$count = 30014;
	#10 counter$count = 30015;
	#10 counter$count = 30016;
	#10 counter$count = 30017;
	#10 counter$count = 30018;
	#10 counter$count = 30019;
	#10 counter$count = 30020;
	#10 counter$count = 30021;
	#10 counter$count = 30022;
	#10 counter$count = 30023;
	#10 counter$count = 30024;
	#10 counter$count = 30025;
	#10 counter$count = 30026;
	#10 counter$count = 30027;
	#10 counter$count = 30028;
	#10 counter$count = 30029;
	#10 counter$count = 30030;
	#10 counter$count = 30031;
	#10 counter$count = 30032;
	#10 counter$count = 30033;
	#10 counter$count = 30034;
	#10 counter$count = 30035;
	#10 counter$count = 30036;
	#10 counter$count = 30037;
	#10 counter$count = 30038;
	#10 counter$count = 30039;
	#10 counter$count = 30040;
	#10 counter$count = 30041;
	#10 counter$count = 30042;
	#10 counter$count = 30043;
	#10 counter$count = 30044;
	#10 counter$count = 30045;
	#10 counter$count = 30046;
	#10 counter$count = 30047;
	#10 counter$count = 30048;
	#10 counter$count = 30049;
	#10 counter$count = 30050;
	#10 counter$count = 30051;
	#10 counter$count = 30052;
	#10 counter$count = 30053;
	#10 counter$count = 30054;
	#10 counter$count = 30055;
	#10 counter$count = 30056;
	#10 counter$count = 30057;
	#10 counter$count = 30058;
	#10 counter$count = 30059;
	#10 counter$count = 30060;
	#10 counter$count = 30061;
	#10 counter$count = 30062;
	#10 counter$count = 30063;
	#10 counter$count = 30064;
	#10 counter$count = 30065;
	#10 counter$count = 30066;
	#10 counter$count = 30067;
	#10 counter$count = 30068;
	#10 counter$count = 30069;
	#10 counter$count = 30070;
	#10 counter$count = 30071;
	#10 counter$count = 30072;
	#10 counter$count = 30073;
	#10 counter$count = 30074;
	#10 counter$count = 30075;
	#10 counter$count = 30076;
	#10 counter$count = 30077;
	#10 counter$count = 30078;
	#10 counter$count = 30079;
	#10 counter$count = 30080;
	#10 counter$count = 30081;
	#10 counter$count = 30082;
	#10 counter$count = 30083;
	#10 counter$count = 30084;
	#10 counter$count = 30085;
	#10 counter$count = 30086;
	#10 counter$count = 30087;
	#10 counter$count = 30088;
	#10 counter$count = 30089;
	#10 counter$count = 30090;
	#10 counter$count = 30091;
	#10 counter$count = 30092;
	#10 counter$count = 30093;
	#10 counter$count = 30094;
	#10 counter$count = 30095;
	#10 counter$count = 30096;
	#10 counter$count = 30097;
	#10 counter$count = 30098;
	#10 counter$count = 30099;
	#10 counter$count = 30100;
	#10 counter$count = 30101;
	#10 counter$count = 30102;
	#10 counter$count = 30103;
	#10 counter$count = 30104;
	#10 counter$count = 30105;
	#10 counter$count = 30106;
	#10 counter$count = 30107;
	#10 counter$count = 30108;
	#10 counter$count = 30109;
	#10 counter$count = 30110;
	#10 counter$count = 30111;
	#10 counter$count = 30112;
	#10 counter$count = 30113;
	#10 counter$count = 30114;
	#10 counter$count = 30115;
	#10 counter$count = 30116;
	#10 counter$count = 30117;
	#10 counter$count = 30118;
	#10 counter$count = 30119;
	#10 counter$count = 30120;
	#10 counter$count = 30121;
	#10 counter$count = 30122;
	#10 counter$count = 30123;
	#10 counter$count = 30124;
	#10 counter$count = 30125;
	#10 counter$count = 30126;
	#10 counter$count = 30127;
	#10 counter$count = 30128;
	#10 counter$count = 30129;
	#10 counter$count = 30130;
	#10 counter$count = 30131;
	#10 counter$count = 30132;
	#10 counter$count = 30133;
	#10 counter$count = 30134;
	#10 counter$count = 30135;
	#10 counter$count = 30136;
	#10 counter$count = 30137;
	#10 counter$count = 30138;
	#10 counter$count = 30139;
	#10 counter$count = 30140;
	#10 counter$count = 30141;
	#10 counter$count = 30142;
	#10 counter$count = 30143;
	#10 counter$count = 30144;
	#10 counter$count = 30145;
	#10 counter$count = 30146;
	#10 counter$count = 30147;
	#10 counter$count = 30148;
	#10 counter$count = 30149;
	#10 counter$count = 30150;
	#10 counter$count = 30151;
	#10 counter$count = 30152;
	#10 counter$count = 30153;
	#10 counter$count = 30154;
	#10 counter$count = 30155;
	#10 counter$count = 30156;
	#10 counter$count = 30157;
	#10 counter$count = 30158;
	#10 counter$count = 30159;
	#10 counter$count = 30160;
	#10 counter$count = 30161;
	#10 counter$count = 30162;
	#10 counter$count = 30163;
	#10 counter$count = 30164;
	#10 counter$count = 30165;
	#10 counter$count = 30166;
	#10 counter$count = 30167;
	#10 counter$count = 30168;
	#10 counter$count = 30169;
	#10 counter$count = 30170;
	#10 counter$count = 30171;
	#10 counter$count = 30172;
	#10 counter$count = 30173;
	#10 counter$count = 30174;
	#10 counter$count = 30175;
	#10 counter$count = 30176;
	#10 counter$count = 30177;
	#10 counter$count = 30178;
	#10 counter$count = 30179;
	#10 counter$count = 30180;
	#10 counter$count = 30181;
	#10 counter$count = 30182;
	#10 counter$count = 30183;
	#10 counter$count = 30184;
	#10 counter$count = 30185;
	#10 counter$count = 30186;
	#10 counter$count = 30187;
	#10 counter$count = 30188;
	#10 counter$count = 30189;
	#10 counter$count = 30190;
	#10 counter$count = 30191;
	#10 counter$count = 30192;
	#10 counter$count = 30193;
	#10 counter$count = 30194;
	#10 counter$count = 30195;
	#10 counter$count = 30196;
	#10 counter$count = 30197;
	#10 counter$count = 30198;
	#10 counter$count = 30199;
	#10 counter$count = 30200;
	#10 counter$count = 30201;
	#10 counter$count = 30202;
	#10 counter$count = 30203;
	#10 counter$count = 30204;
	#10 counter$count = 30205;
	#10 counter$count = 30206;
	#10 counter$count = 30207;
	#10 counter$count = 30208;
	#10 counter$count = 30209;
	#10 counter$count = 30210;
	#10 counter$count = 30211;
	#10 counter$count = 30212;
	#10 counter$count = 30213;
	#10 counter$count = 30214;
	#10 counter$count = 30215;
	#10 counter$count = 30216;
	#10 counter$count = 30217;
	#10 counter$count = 30218;
	#10 counter$count = 30219;
	#10 counter$count = 30220;
	#10 counter$count = 30221;
	#10 counter$count = 30222;
	#10 counter$count = 30223;
	#10 counter$count = 30224;
	#10 counter$count = 30225;
	#10 counter$count = 30226;
	#10 counter$count = 30227;
	#10 counter$count = 30228;
	#10 counter$count = 30229;
	#10 counter$count = 30230;
	#10 counter$count = 30231;
	#10 counter$count = 30232;
	#10 counter$count = 30233;
	#10 counter$count = 30234;
	#10 counter$count = 30235;
	#10 counter$count = 30236;
	#10 counter$count = 30237;
	#10 counter$count = 30238;
	#10 counter$count = 30239;
	#10 counter$count = 30240;
	#10 counter$count = 30241;
	#10 counter$count = 30242;
	#10 counter$count = 30243;
	#10 counter$count = 30244;
	#10 counter$count = 30245;
	#10 counter$count = 30246;
	#10 counter$count = 30247;
	#10 counter$count = 30248;
	#10 counter$count = 30249;
	#10 counter$count = 30250;
	#10 counter$count = 30251;
	#10 counter$count = 30252;
	#10 counter$count = 30253;
	#10 counter$count = 30254;
	#10 counter$count = 30255;
	#10 counter$count = 30256;
	#10 counter$count = 30257;
	#10 counter$count = 30258;
	#10 counter$count = 30259;
	#10 counter$count = 30260;
	#10 counter$count = 30261;
	#10 counter$count = 30262;
	#10 counter$count = 30263;
	#10 counter$count = 30264;
	#10 counter$count = 30265;
	#10 counter$count = 30266;
	#10 counter$count = 30267;
	#10 counter$count = 30268;
	#10 counter$count = 30269;
	#10 counter$count = 30270;
	#10 counter$count = 30271;
	#10 counter$count = 30272;
	#10 counter$count = 30273;
	#10 counter$count = 30274;
	#10 counter$count = 30275;
	#10 counter$count = 30276;
	#10 counter$count = 30277;
	#10 counter$count = 30278;
	#10 counter$count = 30279;
	#10 counter$count = 30280;
	#10 counter$count = 30281;
	#10 counter$count = 30282;
	#10 counter$count = 30283;
	#10 counter$count = 30284;
	#10 counter$count = 30285;
	#10 counter$count = 30286;
	#10 counter$count = 30287;
	#10 counter$count = 30288;
	#10 counter$count = 30289;
	#10 counter$count = 30290;
	#10 counter$count = 30291;
	#10 counter$count = 30292;
	#10 counter$count = 30293;
	#10 counter$count = 30294;
	#10 counter$count = 30295;
	#10 counter$count = 30296;
	#10 counter$count = 30297;
	#10 counter$count = 30298;
	#10 counter$count = 30299;
	#10 counter$count = 30300;
	#10 counter$count = 30301;
	#10 counter$count = 30302;
	#10 counter$count = 30303;
	#10 counter$count = 30304;
	#10 counter$count = 30305;
	#10 counter$count = 30306;
	#10 counter$count = 30307;
	#10 counter$count = 30308;
	#10 counter$count = 30309;
	#10 counter$count = 30310;
	#10 counter$count = 30311;
	#10 counter$count = 30312;
	#10 counter$count = 30313;
	#10 counter$count = 30314;
	#10 counter$count = 30315;
	#10 counter$count = 30316;
	#10 counter$count = 30317;
	#10 counter$count = 30318;
	#10 counter$count = 30319;
	#10 counter$count = 30320;
	#10 counter$count = 30321;
	#10 counter$count = 30322;
	#10 counter$count = 30323;
	#10 counter$count = 30324;
	#10 counter$count = 30325;
	#10 counter$count = 30326;
	#10 counter$count = 30327;
	#10 counter$count = 30328;
	#10 counter$count = 30329;
	#10 counter$count = 30330;
	#10 counter$count = 30331;
	#10 counter$count = 30332;
	#10 counter$count = 30333;
	#10 counter$count = 30334;
	#10 counter$count = 30335;
	#10 counter$count = 30336;
	#10 counter$count = 30337;
	#10 counter$count = 30338;
	#10 counter$count = 30339;
	#10 counter$count = 30340;
	#10 counter$count = 30341;
	#10 counter$count = 30342;
	#10 counter$count = 30343;
	#10 counter$count = 30344;
	#10 counter$count = 30345;
	#10 counter$count = 30346;
	#10 counter$count = 30347;
	#10 counter$count = 30348;
	#10 counter$count = 30349;
	#10 counter$count = 30350;
	#10 counter$count = 30351;
	#10 counter$count = 30352;
	#10 counter$count = 30353;
	#10 counter$count = 30354;
	#10 counter$count = 30355;
	#10 counter$count = 30356;
	#10 counter$count = 30357;
	#10 counter$count = 30358;
	#10 counter$count = 30359;
	#10 counter$count = 30360;
	#10 counter$count = 30361;
	#10 counter$count = 30362;
	#10 counter$count = 30363;
	#10 counter$count = 30364;
	#10 counter$count = 30365;
	#10 counter$count = 30366;
	#10 counter$count = 30367;
	#10 counter$count = 30368;
	#10 counter$count = 30369;
	#10 counter$count = 30370;
	#10 counter$count = 30371;
	#10 counter$count = 30372;
	#10 counter$count = 30373;
	#10 counter$count = 30374;
	#10 counter$count = 30375;
	#10 counter$count = 30376;
	#10 counter$count = 30377;
	#10 counter$count = 30378;
	#10 counter$count = 30379;
	#10 counter$count = 30380;
	#10 counter$count = 30381;
	#10 counter$count = 30382;
	#10 counter$count = 30383;
	#10 counter$count = 30384;
	#10 counter$count = 30385;
	#10 counter$count = 30386;
	#10 counter$count = 30387;
	#10 counter$count = 30388;
	#10 counter$count = 30389;
	#10 counter$count = 30390;
	#10 counter$count = 30391;
	#10 counter$count = 30392;
	#10 counter$count = 30393;
	#10 counter$count = 30394;
	#10 counter$count = 30395;
	#10 counter$count = 30396;
	#10 counter$count = 30397;
	#10 counter$count = 30398;
	#10 counter$count = 30399;
	#10 counter$count = 30400;
	#10 counter$count = 30401;
	#10 counter$count = 30402;
	#10 counter$count = 30403;
	#10 counter$count = 30404;
	#10 counter$count = 30405;
	#10 counter$count = 30406;
	#10 counter$count = 30407;
	#10 counter$count = 30408;
	#10 counter$count = 30409;
	#10 counter$count = 30410;
	#10 counter$count = 30411;
	#10 counter$count = 30412;
	#10 counter$count = 30413;
	#10 counter$count = 30414;
	#10 counter$count = 30415;
	#10 counter$count = 30416;
	#10 counter$count = 30417;
	#10 counter$count = 30418;
	#10 counter$count = 30419;
	#10 counter$count = 30420;
	#10 counter$count = 30421;
	#10 counter$count = 30422;
	#10 counter$count = 30423;
	#10 counter$count = 30424;
	#10 counter$count = 30425;
	#10 counter$count = 30426;
	#10 counter$count = 30427;
	#10 counter$count = 30428;
	#10 counter$count = 30429;
	#10 counter$count = 30430;
	#10 counter$count = 30431;
	#10 counter$count = 30432;
	#10 counter$count = 30433;
	#10 counter$count = 30434;
	#10 counter$count = 30435;
	#10 counter$count = 30436;
	#10 counter$count = 30437;
	#10 counter$count = 30438;
	#10 counter$count = 30439;
	#10 counter$count = 30440;
	#10 counter$count = 30441;
	#10 counter$count = 30442;
	#10 counter$count = 30443;
	#10 counter$count = 30444;
	#10 counter$count = 30445;
	#10 counter$count = 30446;
	#10 counter$count = 30447;
	#10 counter$count = 30448;
	#10 counter$count = 30449;
	#10 counter$count = 30450;
	#10 counter$count = 30451;
	#10 counter$count = 30452;
	#10 counter$count = 30453;
	#10 counter$count = 30454;
	#10 counter$count = 30455;
	#10 counter$count = 30456;
	#10 counter$count = 30457;
	#10 counter$count = 30458;
	#10 counter$count = 30459;
	#10 counter$count = 30460;
	#10 counter$count = 30461;
	#10 counter$count = 30462;
	#10 counter$count = 30463;
	#10 counter$count = 30464;
	#10 counter$count = 30465;
	#10 counter$count = 30466;
	#10 counter$count = 30467;
	#10 counter$count = 30468;
	#10 counter$count = 30469;
	#10 counter$count = 30470;
	#10 counter$count = 30471;
	#10 counter$count = 30472;
	#10 counter$count = 30473;
	#10 counter$count = 30474;
	#10 counter$count = 30475;
	#10 counter$count = 30476;
	#10 counter$count = 30477;
	#10 counter$count = 30478;
	#10 counter$count = 30479;
	#10 counter$count = 30480;
	#10 counter$count = 30481;
	#10 counter$count = 30482;
	#10 counter$count = 30483;
	#10 counter$count = 30484;
	#10 counter$count = 30485;
	#10 counter$count = 30486;
	#10 counter$count = 30487;
	#10 counter$count = 30488;
	#10 counter$count = 30489;
	#10 counter$count = 30490;
	#10 counter$count = 30491;
	#10 counter$count = 30492;
	#10 counter$count = 30493;
	#10 counter$count = 30494;
	#10 counter$count = 30495;
	#10 counter$count = 30496;
	#10 counter$count = 30497;
	#10 counter$count = 30498;
	#10 counter$count = 30499;
	#10 counter$count = 30500;
	#10 counter$count = 30501;
	#10 counter$count = 30502;
	#10 counter$count = 30503;
	#10 counter$count = 30504;
	#10 counter$count = 30505;
	#10 counter$count = 30506;
	#10 counter$count = 30507;
	#10 counter$count = 30508;
	#10 counter$count = 30509;
	#10 counter$count = 30510;
	#10 counter$count = 30511;
	#10 counter$count = 30512;
	#10 counter$count = 30513;
	#10 counter$count = 30514;
	#10 counter$count = 30515;
	#10 counter$count = 30516;
	#10 counter$count = 30517;
	#10 counter$count = 30518;
	#10 counter$count = 30519;
	#10 counter$count = 30520;
	#10 counter$count = 30521;
	#10 counter$count = 30522;
	#10 counter$count = 30523;
	#10 counter$count = 30524;
	#10 counter$count = 30525;
	#10 counter$count = 30526;
	#10 counter$count = 30527;
	#10 counter$count = 30528;
	#10 counter$count = 30529;
	#10 counter$count = 30530;
	#10 counter$count = 30531;
	#10 counter$count = 30532;
	#10 counter$count = 30533;
	#10 counter$count = 30534;
	#10 counter$count = 30535;
	#10 counter$count = 30536;
	#10 counter$count = 30537;
	#10 counter$count = 30538;
	#10 counter$count = 30539;
	#10 counter$count = 30540;
	#10 counter$count = 30541;
	#10 counter$count = 30542;
	#10 counter$count = 30543;
	#10 counter$count = 30544;
	#10 counter$count = 30545;
	#10 counter$count = 30546;
	#10 counter$count = 30547;
	#10 counter$count = 30548;
	#10 counter$count = 30549;
	#10 counter$count = 30550;
	#10 counter$count = 30551;
	#10 counter$count = 30552;
	#10 counter$count = 30553;
	#10 counter$count = 30554;
	#10 counter$count = 30555;
	#10 counter$count = 30556;
	#10 counter$count = 30557;
	#10 counter$count = 30558;
	#10 counter$count = 30559;
	#10 counter$count = 30560;
	#10 counter$count = 30561;
	#10 counter$count = 30562;
	#10 counter$count = 30563;
	#10 counter$count = 30564;
	#10 counter$count = 30565;
	#10 counter$count = 30566;
	#10 counter$count = 30567;
	#10 counter$count = 30568;
	#10 counter$count = 30569;
	#10 counter$count = 30570;
	#10 counter$count = 30571;
	#10 counter$count = 30572;
	#10 counter$count = 30573;
	#10 counter$count = 30574;
	#10 counter$count = 30575;
	#10 counter$count = 30576;
	#10 counter$count = 30577;
	#10 counter$count = 30578;
	#10 counter$count = 30579;
	#10 counter$count = 30580;
	#10 counter$count = 30581;
	#10 counter$count = 30582;
	#10 counter$count = 30583;
	#10 counter$count = 30584;
	#10 counter$count = 30585;
	#10 counter$count = 30586;
	#10 counter$count = 30587;
	#10 counter$count = 30588;
	#10 counter$count = 30589;
	#10 counter$count = 30590;
	#10 counter$count = 30591;
	#10 counter$count = 30592;
	#10 counter$count = 30593;
	#10 counter$count = 30594;
	#10 counter$count = 30595;
	#10 counter$count = 30596;
	#10 counter$count = 30597;
	#10 counter$count = 30598;
	#10 counter$count = 30599;
	#10 counter$count = 30600;
	#10 counter$count = 30601;
	#10 counter$count = 30602;
	#10 counter$count = 30603;
	#10 counter$count = 30604;
	#10 counter$count = 30605;
	#10 counter$count = 30606;
	#10 counter$count = 30607;
	#10 counter$count = 30608;
	#10 counter$count = 30609;
	#10 counter$count = 30610;
	#10 counter$count = 30611;
	#10 counter$count = 30612;
	#10 counter$count = 30613;
	#10 counter$count = 30614;
	#10 counter$count = 30615;
	#10 counter$count = 30616;
	#10 counter$count = 30617;
	#10 counter$count = 30618;
	#10 counter$count = 30619;
	#10 counter$count = 30620;
	#10 counter$count = 30621;
	#10 counter$count = 30622;
	#10 counter$count = 30623;
	#10 counter$count = 30624;
	#10 counter$count = 30625;
	#10 counter$count = 30626;
	#10 counter$count = 30627;
	#10 counter$count = 30628;
	#10 counter$count = 30629;
	#10 counter$count = 30630;
	#10 counter$count = 30631;
	#10 counter$count = 30632;
	#10 counter$count = 30633;
	#10 counter$count = 30634;
	#10 counter$count = 30635;
	#10 counter$count = 30636;
	#10 counter$count = 30637;
	#10 counter$count = 30638;
	#10 counter$count = 30639;
	#10 counter$count = 30640;
	#10 counter$count = 30641;
	#10 counter$count = 30642;
	#10 counter$count = 30643;
	#10 counter$count = 30644;
	#10 counter$count = 30645;
	#10 counter$count = 30646;
	#10 counter$count = 30647;
	#10 counter$count = 30648;
	#10 counter$count = 30649;
	#10 counter$count = 30650;
	#10 counter$count = 30651;
	#10 counter$count = 30652;
	#10 counter$count = 30653;
	#10 counter$count = 30654;
	#10 counter$count = 30655;
	#10 counter$count = 30656;
	#10 counter$count = 30657;
	#10 counter$count = 30658;
	#10 counter$count = 30659;
	#10 counter$count = 30660;
	#10 counter$count = 30661;
	#10 counter$count = 30662;
	#10 counter$count = 30663;
	#10 counter$count = 30664;
	#10 counter$count = 30665;
	#10 counter$count = 30666;
	#10 counter$count = 30667;
	#10 counter$count = 30668;
	#10 counter$count = 30669;
	#10 counter$count = 30670;
	#10 counter$count = 30671;
	#10 counter$count = 30672;
	#10 counter$count = 30673;
	#10 counter$count = 30674;
	#10 counter$count = 30675;
	#10 counter$count = 30676;
	#10 counter$count = 30677;
	#10 counter$count = 30678;
	#10 counter$count = 30679;
	#10 counter$count = 30680;
	#10 counter$count = 30681;
	#10 counter$count = 30682;
	#10 counter$count = 30683;
	#10 counter$count = 30684;
	#10 counter$count = 30685;
	#10 counter$count = 30686;
	#10 counter$count = 30687;
	#10 counter$count = 30688;
	#10 counter$count = 30689;
	#10 counter$count = 30690;
	#10 counter$count = 30691;
	#10 counter$count = 30692;
	#10 counter$count = 30693;
	#10 counter$count = 30694;
	#10 counter$count = 30695;
	#10 counter$count = 30696;
	#10 counter$count = 30697;
	#10 counter$count = 30698;
	#10 counter$count = 30699;
	#10 counter$count = 30700;
	#10 counter$count = 30701;
	#10 counter$count = 30702;
	#10 counter$count = 30703;
	#10 counter$count = 30704;
	#10 counter$count = 30705;
	#10 counter$count = 30706;
	#10 counter$count = 30707;
	#10 counter$count = 30708;
	#10 counter$count = 30709;
	#10 counter$count = 30710;
	#10 counter$count = 30711;
	#10 counter$count = 30712;
	#10 counter$count = 30713;
	#10 counter$count = 30714;
	#10 counter$count = 30715;
	#10 counter$count = 30716;
	#10 counter$count = 30717;
	#10 counter$count = 30718;
	#10 counter$count = 30719;
	#10 counter$count = 30720;
	#10 counter$count = 30721;
	#10 counter$count = 30722;
	#10 counter$count = 30723;
	#10 counter$count = 30724;
	#10 counter$count = 30725;
	#10 counter$count = 30726;
	#10 counter$count = 30727;
	#10 counter$count = 30728;
	#10 counter$count = 30729;
	#10 counter$count = 30730;
	#10 counter$count = 30731;
	#10 counter$count = 30732;
	#10 counter$count = 30733;
	#10 counter$count = 30734;
	#10 counter$count = 30735;
	#10 counter$count = 30736;
	#10 counter$count = 30737;
	#10 counter$count = 30738;
	#10 counter$count = 30739;
	#10 counter$count = 30740;
	#10 counter$count = 30741;
	#10 counter$count = 30742;
	#10 counter$count = 30743;
	#10 counter$count = 30744;
	#10 counter$count = 30745;
	#10 counter$count = 30746;
	#10 counter$count = 30747;
	#10 counter$count = 30748;
	#10 counter$count = 30749;
	#10 counter$count = 30750;
	#10 counter$count = 30751;
	#10 counter$count = 30752;
	#10 counter$count = 30753;
	#10 counter$count = 30754;
	#10 counter$count = 30755;
	#10 counter$count = 30756;
	#10 counter$count = 30757;
	#10 counter$count = 30758;
	#10 counter$count = 30759;
	#10 counter$count = 30760;
	#10 counter$count = 30761;
	#10 counter$count = 30762;
	#10 counter$count = 30763;
	#10 counter$count = 30764;
	#10 counter$count = 30765;
	#10 counter$count = 30766;
	#10 counter$count = 30767;
	#10 counter$count = 30768;
	#10 counter$count = 30769;
	#10 counter$count = 30770;
	#10 counter$count = 30771;
	#10 counter$count = 30772;
	#10 counter$count = 30773;
	#10 counter$count = 30774;
	#10 counter$count = 30775;
	#10 counter$count = 30776;
	#10 counter$count = 30777;
	#10 counter$count = 30778;
	#10 counter$count = 30779;
	#10 counter$count = 30780;
	#10 counter$count = 30781;
	#10 counter$count = 30782;
	#10 counter$count = 30783;
	#10 counter$count = 30784;
	#10 counter$count = 30785;
	#10 counter$count = 30786;
	#10 counter$count = 30787;
	#10 counter$count = 30788;
	#10 counter$count = 30789;
	#10 counter$count = 30790;
	#10 counter$count = 30791;
	#10 counter$count = 30792;
	#10 counter$count = 30793;
	#10 counter$count = 30794;
	#10 counter$count = 30795;
	#10 counter$count = 30796;
	#10 counter$count = 30797;
	#10 counter$count = 30798;
	#10 counter$count = 30799;
	#10 counter$count = 30800;
	#10 counter$count = 30801;
	#10 counter$count = 30802;
	#10 counter$count = 30803;
	#10 counter$count = 30804;
	#10 counter$count = 30805;
	#10 counter$count = 30806;
	#10 counter$count = 30807;
	#10 counter$count = 30808;
	#10 counter$count = 30809;
	#10 counter$count = 30810;
	#10 counter$count = 30811;
	#10 counter$count = 30812;
	#10 counter$count = 30813;
	#10 counter$count = 30814;
	#10 counter$count = 30815;
	#10 counter$count = 30816;
	#10 counter$count = 30817;
	#10 counter$count = 30818;
	#10 counter$count = 30819;
	#10 counter$count = 30820;
	#10 counter$count = 30821;
	#10 counter$count = 30822;
	#10 counter$count = 30823;
	#10 counter$count = 30824;
	#10 counter$count = 30825;
	#10 counter$count = 30826;
	#10 counter$count = 30827;
	#10 counter$count = 30828;
	#10 counter$count = 30829;
	#10 counter$count = 30830;
	#10 counter$count = 30831;
	#10 counter$count = 30832;
	#10 counter$count = 30833;
	#10 counter$count = 30834;
	#10 counter$count = 30835;
	#10 counter$count = 30836;
	#10 counter$count = 30837;
	#10 counter$count = 30838;
	#10 counter$count = 30839;
	#10 counter$count = 30840;
	#10 counter$count = 30841;
	#10 counter$count = 30842;
	#10 counter$count = 30843;
	#10 counter$count = 30844;
	#10 counter$count = 30845;
	#10 counter$count = 30846;
	#10 counter$count = 30847;
	#10 counter$count = 30848;
	#10 counter$count = 30849;
	#10 counter$count = 30850;
	#10 counter$count = 30851;
	#10 counter$count = 30852;
	#10 counter$count = 30853;
	#10 counter$count = 30854;
	#10 counter$count = 30855;
	#10 counter$count = 30856;
	#10 counter$count = 30857;
	#10 counter$count = 30858;
	#10 counter$count = 30859;
	#10 counter$count = 30860;
	#10 counter$count = 30861;
	#10 counter$count = 30862;
	#10 counter$count = 30863;
	#10 counter$count = 30864;
	#10 counter$count = 30865;
	#10 counter$count = 30866;
	#10 counter$count = 30867;
	#10 counter$count = 30868;
	#10 counter$count = 30869;
	#10 counter$count = 30870;
	#10 counter$count = 30871;
	#10 counter$count = 30872;
	#10 counter$count = 30873;
	#10 counter$count = 30874;
	#10 counter$count = 30875;
	#10 counter$count = 30876;
	#10 counter$count = 30877;
	#10 counter$count = 30878;
	#10 counter$count = 30879;
	#10 counter$count = 30880;
	#10 counter$count = 30881;
	#10 counter$count = 30882;
	#10 counter$count = 30883;
	#10 counter$count = 30884;
	#10 counter$count = 30885;
	#10 counter$count = 30886;
	#10 counter$count = 30887;
	#10 counter$count = 30888;
	#10 counter$count = 30889;
	#10 counter$count = 30890;
	#10 counter$count = 30891;
	#10 counter$count = 30892;
	#10 counter$count = 30893;
	#10 counter$count = 30894;
	#10 counter$count = 30895;
	#10 counter$count = 30896;
	#10 counter$count = 30897;
	#10 counter$count = 30898;
	#10 counter$count = 30899;
	#10 counter$count = 30900;
	#10 counter$count = 30901;
	#10 counter$count = 30902;
	#10 counter$count = 30903;
	#10 counter$count = 30904;
	#10 counter$count = 30905;
	#10 counter$count = 30906;
	#10 counter$count = 30907;
	#10 counter$count = 30908;
	#10 counter$count = 30909;
	#10 counter$count = 30910;
	#10 counter$count = 30911;
	#10 counter$count = 30912;
	#10 counter$count = 30913;
	#10 counter$count = 30914;
	#10 counter$count = 30915;
	#10 counter$count = 30916;
	#10 counter$count = 30917;
	#10 counter$count = 30918;
	#10 counter$count = 30919;
	#10 counter$count = 30920;
	#10 counter$count = 30921;
	#10 counter$count = 30922;
	#10 counter$count = 30923;
	#10 counter$count = 30924;
	#10 counter$count = 30925;
	#10 counter$count = 30926;
	#10 counter$count = 30927;
	#10 counter$count = 30928;
	#10 counter$count = 30929;
	#10 counter$count = 30930;
	#10 counter$count = 30931;
	#10 counter$count = 30932;
	#10 counter$count = 30933;
	#10 counter$count = 30934;
	#10 counter$count = 30935;
	#10 counter$count = 30936;
	#10 counter$count = 30937;
	#10 counter$count = 30938;
	#10 counter$count = 30939;
	#10 counter$count = 30940;
	#10 counter$count = 30941;
	#10 counter$count = 30942;
	#10 counter$count = 30943;
	#10 counter$count = 30944;
	#10 counter$count = 30945;
	#10 counter$count = 30946;
	#10 counter$count = 30947;
	#10 counter$count = 30948;
	#10 counter$count = 30949;
	#10 counter$count = 30950;
	#10 counter$count = 30951;
	#10 counter$count = 30952;
	#10 counter$count = 30953;
	#10 counter$count = 30954;
	#10 counter$count = 30955;
	#10 counter$count = 30956;
	#10 counter$count = 30957;
	#10 counter$count = 30958;
	#10 counter$count = 30959;
	#10 counter$count = 30960;
	#10 counter$count = 30961;
	#10 counter$count = 30962;
	#10 counter$count = 30963;
	#10 counter$count = 30964;
	#10 counter$count = 30965;
	#10 counter$count = 30966;
	#10 counter$count = 30967;
	#10 counter$count = 30968;
	#10 counter$count = 30969;
	#10 counter$count = 30970;
	#10 counter$count = 30971;
	#10 counter$count = 30972;
	#10 counter$count = 30973;
	#10 counter$count = 30974;
	#10 counter$count = 30975;
	#10 counter$count = 30976;
	#10 counter$count = 30977;
	#10 counter$count = 30978;
	#10 counter$count = 30979;
	#10 counter$count = 30980;
	#10 counter$count = 30981;
	#10 counter$count = 30982;
	#10 counter$count = 30983;
	#10 counter$count = 30984;
	#10 counter$count = 30985;
	#10 counter$count = 30986;
	#10 counter$count = 30987;
	#10 counter$count = 30988;
	#10 counter$count = 30989;
	#10 counter$count = 30990;
	#10 counter$count = 30991;
	#10 counter$count = 30992;
	#10 counter$count = 30993;
	#10 counter$count = 30994;
	#10 counter$count = 30995;
	#10 counter$count = 30996;
	#10 counter$count = 30997;
	#10 counter$count = 30998;
	#10 counter$count = 30999;
	#10 counter$count = 31000;
	#10 counter$count = 31001;
	#10 counter$count = 31002;
	#10 counter$count = 31003;
	#10 counter$count = 31004;
	#10 counter$count = 31005;
	#10 counter$count = 31006;
	#10 counter$count = 31007;
	#10 counter$count = 31008;
	#10 counter$count = 31009;
	#10 counter$count = 31010;
	#10 counter$count = 31011;
	#10 counter$count = 31012;
	#10 counter$count = 31013;
	#10 counter$count = 31014;
	#10 counter$count = 31015;
	#10 counter$count = 31016;
	#10 counter$count = 31017;
	#10 counter$count = 31018;
	#10 counter$count = 31019;
	#10 counter$count = 31020;
	#10 counter$count = 31021;
	#10 counter$count = 31022;
	#10 counter$count = 31023;
	#10 counter$count = 31024;
	#10 counter$count = 31025;
	#10 counter$count = 31026;
	#10 counter$count = 31027;
	#10 counter$count = 31028;
	#10 counter$count = 31029;
	#10 counter$count = 31030;
	#10 counter$count = 31031;
	#10 counter$count = 31032;
	#10 counter$count = 31033;
	#10 counter$count = 31034;
	#10 counter$count = 31035;
	#10 counter$count = 31036;
	#10 counter$count = 31037;
	#10 counter$count = 31038;
	#10 counter$count = 31039;
	#10 counter$count = 31040;
	#10 counter$count = 31041;
	#10 counter$count = 31042;
	#10 counter$count = 31043;
	#10 counter$count = 31044;
	#10 counter$count = 31045;
	#10 counter$count = 31046;
	#10 counter$count = 31047;
	#10 counter$count = 31048;
	#10 counter$count = 31049;
	#10 counter$count = 31050;
	#10 counter$count = 31051;
	#10 counter$count = 31052;
	#10 counter$count = 31053;
	#10 counter$count = 31054;
	#10 counter$count = 31055;
	#10 counter$count = 31056;
	#10 counter$count = 31057;
	#10 counter$count = 31058;
	#10 counter$count = 31059;
	#10 counter$count = 31060;
	#10 counter$count = 31061;
	#10 counter$count = 31062;
	#10 counter$count = 31063;
	#10 counter$count = 31064;
	#10 counter$count = 31065;
	#10 counter$count = 31066;
	#10 counter$count = 31067;
	#10 counter$count = 31068;
	#10 counter$count = 31069;
	#10 counter$count = 31070;
	#10 counter$count = 31071;
	#10 counter$count = 31072;
	#10 counter$count = 31073;
	#10 counter$count = 31074;
	#10 counter$count = 31075;
	#10 counter$count = 31076;
	#10 counter$count = 31077;
	#10 counter$count = 31078;
	#10 counter$count = 31079;
	#10 counter$count = 31080;
	#10 counter$count = 31081;
	#10 counter$count = 31082;
	#10 counter$count = 31083;
	#10 counter$count = 31084;
	#10 counter$count = 31085;
	#10 counter$count = 31086;
	#10 counter$count = 31087;
	#10 counter$count = 31088;
	#10 counter$count = 31089;
	#10 counter$count = 31090;
	#10 counter$count = 31091;
	#10 counter$count = 31092;
	#10 counter$count = 31093;
	#10 counter$count = 31094;
	#10 counter$count = 31095;
	#10 counter$count = 31096;
	#10 counter$count = 31097;
	#10 counter$count = 31098;
	#10 counter$count = 31099;
	#10 counter$count = 31100;
	#10 counter$count = 31101;
	#10 counter$count = 31102;
	#10 counter$count = 31103;
	#10 counter$count = 31104;
	#10 counter$count = 31105;
	#10 counter$count = 31106;
	#10 counter$count = 31107;
	#10 counter$count = 31108;
	#10 counter$count = 31109;
	#10 counter$count = 31110;
	#10 counter$count = 31111;
	#10 counter$count = 31112;
	#10 counter$count = 31113;
	#10 counter$count = 31114;
	#10 counter$count = 31115;
	#10 counter$count = 31116;
	#10 counter$count = 31117;
	#10 counter$count = 31118;
	#10 counter$count = 31119;
	#10 counter$count = 31120;
	#10 counter$count = 31121;
	#10 counter$count = 31122;
	#10 counter$count = 31123;
	#10 counter$count = 31124;
	#10 counter$count = 31125;
	#10 counter$count = 31126;
	#10 counter$count = 31127;
	#10 counter$count = 31128;
	#10 counter$count = 31129;
	#10 counter$count = 31130;
	#10 counter$count = 31131;
	#10 counter$count = 31132;
	#10 counter$count = 31133;
	#10 counter$count = 31134;
	#10 counter$count = 31135;
	#10 counter$count = 31136;
	#10 counter$count = 31137;
	#10 counter$count = 31138;
	#10 counter$count = 31139;
	#10 counter$count = 31140;
	#10 counter$count = 31141;
	#10 counter$count = 31142;
	#10 counter$count = 31143;
	#10 counter$count = 31144;
	#10 counter$count = 31145;
	#10 counter$count = 31146;
	#10 counter$count = 31147;
	#10 counter$count = 31148;
	#10 counter$count = 31149;
	#10 counter$count = 31150;
	#10 counter$count = 31151;
	#10 counter$count = 31152;
	#10 counter$count = 31153;
	#10 counter$count = 31154;
	#10 counter$count = 31155;
	#10 counter$count = 31156;
	#10 counter$count = 31157;
	#10 counter$count = 31158;
	#10 counter$count = 31159;
	#10 counter$count = 31160;
	#10 counter$count = 31161;
	#10 counter$count = 31162;
	#10 counter$count = 31163;
	#10 counter$count = 31164;
	#10 counter$count = 31165;
	#10 counter$count = 31166;
	#10 counter$count = 31167;
	#10 counter$count = 31168;
	#10 counter$count = 31169;
	#10 counter$count = 31170;
	#10 counter$count = 31171;
	#10 counter$count = 31172;
	#10 counter$count = 31173;
	#10 counter$count = 31174;
	#10 counter$count = 31175;
	#10 counter$count = 31176;
	#10 counter$count = 31177;
	#10 counter$count = 31178;
	#10 counter$count = 31179;
	#10 counter$count = 31180;
	#10 counter$count = 31181;
	#10 counter$count = 31182;
	#10 counter$count = 31183;
	#10 counter$count = 31184;
	#10 counter$count = 31185;
	#10 counter$count = 31186;
	#10 counter$count = 31187;
	#10 counter$count = 31188;
	#10 counter$count = 31189;
	#10 counter$count = 31190;
	#10 counter$count = 31191;
	#10 counter$count = 31192;
	#10 counter$count = 31193;
	#10 counter$count = 31194;
	#10 counter$count = 31195;
	#10 counter$count = 31196;
	#10 counter$count = 31197;
	#10 counter$count = 31198;
	#10 counter$count = 31199;
	#10 counter$count = 31200;
	#10 counter$count = 31201;
	#10 counter$count = 31202;
	#10 counter$count = 31203;
	#10 counter$count = 31204;
	#10 counter$count = 31205;
	#10 counter$count = 31206;
	#10 counter$count = 31207;
	#10 counter$count = 31208;
	#10 counter$count = 31209;
	#10 counter$count = 31210;
	#10 counter$count = 31211;
	#10 counter$count = 31212;
	#10 counter$count = 31213;
	#10 counter$count = 31214;
	#10 counter$count = 31215;
	#10 counter$count = 31216;
	#10 counter$count = 31217;
	#10 counter$count = 31218;
	#10 counter$count = 31219;
	#10 counter$count = 31220;
	#10 counter$count = 31221;
	#10 counter$count = 31222;
	#10 counter$count = 31223;
	#10 counter$count = 31224;
	#10 counter$count = 31225;
	#10 counter$count = 31226;
	#10 counter$count = 31227;
	#10 counter$count = 31228;
	#10 counter$count = 31229;
	#10 counter$count = 31230;
	#10 counter$count = 31231;
	#10 counter$count = 31232;
	#10 counter$count = 31233;
	#10 counter$count = 31234;
	#10 counter$count = 31235;
	#10 counter$count = 31236;
	#10 counter$count = 31237;
	#10 counter$count = 31238;
	#10 counter$count = 31239;
	#10 counter$count = 31240;
	#10 counter$count = 31241;
	#10 counter$count = 31242;
	#10 counter$count = 31243;
	#10 counter$count = 31244;
	#10 counter$count = 31245;
	#10 counter$count = 31246;
	#10 counter$count = 31247;
	#10 counter$count = 31248;
	#10 counter$count = 31249;
	#10 counter$count = 31250;
	#10 counter$count = 31251;
	#10 counter$count = 31252;
	#10 counter$count = 31253;
	#10 counter$count = 31254;
	#10 counter$count = 31255;
	#10 counter$count = 31256;
	#10 counter$count = 31257;
	#10 counter$count = 31258;
	#10 counter$count = 31259;
	#10 counter$count = 31260;
	#10 counter$count = 31261;
	#10 counter$count = 31262;
	#10 counter$count = 31263;
	#10 counter$count = 31264;
	#10 counter$count = 31265;
	#10 counter$count = 31266;
	#10 counter$count = 31267;
	#10 counter$count = 31268;
	#10 counter$count = 31269;
	#10 counter$count = 31270;
	#10 counter$count = 31271;
	#10 counter$count = 31272;
	#10 counter$count = 31273;
	#10 counter$count = 31274;
	#10 counter$count = 31275;
	#10 counter$count = 31276;
	#10 counter$count = 31277;
	#10 counter$count = 31278;
	#10 counter$count = 31279;
	#10 counter$count = 31280;
	#10 counter$count = 31281;
	#10 counter$count = 31282;
	#10 counter$count = 31283;
	#10 counter$count = 31284;
	#10 counter$count = 31285;
	#10 counter$count = 31286;
	#10 counter$count = 31287;
	#10 counter$count = 31288;
	#10 counter$count = 31289;
	#10 counter$count = 31290;
	#10 counter$count = 31291;
	#10 counter$count = 31292;
	#10 counter$count = 31293;
	#10 counter$count = 31294;
	#10 counter$count = 31295;
	#10 counter$count = 31296;
	#10 counter$count = 31297;
	#10 counter$count = 31298;
	#10 counter$count = 31299;
	#10 counter$count = 31300;
	#10 counter$count = 31301;
	#10 counter$count = 31302;
	#10 counter$count = 31303;
	#10 counter$count = 31304;
	#10 counter$count = 31305;
	#10 counter$count = 31306;
	#10 counter$count = 31307;
	#10 counter$count = 31308;
	#10 counter$count = 31309;
	#10 counter$count = 31310;
	#10 counter$count = 31311;
	#10 counter$count = 31312;
	#10 counter$count = 31313;
	#10 counter$count = 31314;
	#10 counter$count = 31315;
	#10 counter$count = 31316;
	#10 counter$count = 31317;
	#10 counter$count = 31318;
	#10 counter$count = 31319;
	#10 counter$count = 31320;
	#10 counter$count = 31321;
	#10 counter$count = 31322;
	#10 counter$count = 31323;
	#10 counter$count = 31324;
	#10 counter$count = 31325;
	#10 counter$count = 31326;
	#10 counter$count = 31327;
	#10 counter$count = 31328;
	#10 counter$count = 31329;
	#10 counter$count = 31330;
	#10 counter$count = 31331;
	#10 counter$count = 31332;
	#10 counter$count = 31333;
	#10 counter$count = 31334;
	#10 counter$count = 31335;
	#10 counter$count = 31336;
	#10 counter$count = 31337;
	#10 counter$count = 31338;
	#10 counter$count = 31339;
	#10 counter$count = 31340;
	#10 counter$count = 31341;
	#10 counter$count = 31342;
	#10 counter$count = 31343;
	#10 counter$count = 31344;
	#10 counter$count = 31345;
	#10 counter$count = 31346;
	#10 counter$count = 31347;
	#10 counter$count = 31348;
	#10 counter$count = 31349;
	#10 counter$count = 31350;
	#10 counter$count = 31351;
	#10 counter$count = 31352;
	#10 counter$count = 31353;
	#10 counter$count = 31354;
	#10 counter$count = 31355;
	#10 counter$count = 31356;
	#10 counter$count = 31357;
	#10 counter$count = 31358;
	#10 counter$count = 31359;
	#10 counter$count = 31360;
	#10 counter$count = 31361;
	#10 counter$count = 31362;
	#10 counter$count = 31363;
	#10 counter$count = 31364;
	#10 counter$count = 31365;
	#10 counter$count = 31366;
	#10 counter$count = 31367;
	#10 counter$count = 31368;
	#10 counter$count = 31369;
	#10 counter$count = 31370;
	#10 counter$count = 31371;
	#10 counter$count = 31372;
	#10 counter$count = 31373;
	#10 counter$count = 31374;
	#10 counter$count = 31375;
	#10 counter$count = 31376;
	#10 counter$count = 31377;
	#10 counter$count = 31378;
	#10 counter$count = 31379;
	#10 counter$count = 31380;
	#10 counter$count = 31381;
	#10 counter$count = 31382;
	#10 counter$count = 31383;
	#10 counter$count = 31384;
	#10 counter$count = 31385;
	#10 counter$count = 31386;
	#10 counter$count = 31387;
	#10 counter$count = 31388;
	#10 counter$count = 31389;
	#10 counter$count = 31390;
	#10 counter$count = 31391;
	#10 counter$count = 31392;
	#10 counter$count = 31393;
	#10 counter$count = 31394;
	#10 counter$count = 31395;
	#10 counter$count = 31396;
	#10 counter$count = 31397;
	#10 counter$count = 31398;
	#10 counter$count = 31399;
	#10 counter$count = 31400;
	#10 counter$count = 31401;
	#10 counter$count = 31402;
	#10 counter$count = 31403;
	#10 counter$count = 31404;
	#10 counter$count = 31405;
	#10 counter$count = 31406;
	#10 counter$count = 31407;
	#10 counter$count = 31408;
	#10 counter$count = 31409;
	#10 counter$count = 31410;
	#10 counter$count = 31411;
	#10 counter$count = 31412;
	#10 counter$count = 31413;
	#10 counter$count = 31414;
	#10 counter$count = 31415;
	#10 counter$count = 31416;
	#10 counter$count = 31417;
	#10 counter$count = 31418;
	#10 counter$count = 31419;
	#10 counter$count = 31420;
	#10 counter$count = 31421;
	#10 counter$count = 31422;
	#10 counter$count = 31423;
	#10 counter$count = 31424;
	#10 counter$count = 31425;
	#10 counter$count = 31426;
	#10 counter$count = 31427;
	#10 counter$count = 31428;
	#10 counter$count = 31429;
	#10 counter$count = 31430;
	#10 counter$count = 31431;
	#10 counter$count = 31432;
	#10 counter$count = 31433;
	#10 counter$count = 31434;
	#10 counter$count = 31435;
	#10 counter$count = 31436;
	#10 counter$count = 31437;
	#10 counter$count = 31438;
	#10 counter$count = 31439;
	#10 counter$count = 31440;
	#10 counter$count = 31441;
	#10 counter$count = 31442;
	#10 counter$count = 31443;
	#10 counter$count = 31444;
	#10 counter$count = 31445;
	#10 counter$count = 31446;
	#10 counter$count = 31447;
	#10 counter$count = 31448;
	#10 counter$count = 31449;
	#10 counter$count = 31450;
	#10 counter$count = 31451;
	#10 counter$count = 31452;
	#10 counter$count = 31453;
	#10 counter$count = 31454;
	#10 counter$count = 31455;
	#10 counter$count = 31456;
	#10 counter$count = 31457;
	#10 counter$count = 31458;
	#10 counter$count = 31459;
	#10 counter$count = 31460;
	#10 counter$count = 31461;
	#10 counter$count = 31462;
	#10 counter$count = 31463;
	#10 counter$count = 31464;
	#10 counter$count = 31465;
	#10 counter$count = 31466;
	#10 counter$count = 31467;
	#10 counter$count = 31468;
	#10 counter$count = 31469;
	#10 counter$count = 31470;
	#10 counter$count = 31471;
	#10 counter$count = 31472;
	#10 counter$count = 31473;
	#10 counter$count = 31474;
	#10 counter$count = 31475;
	#10 counter$count = 31476;
	#10 counter$count = 31477;
	#10 counter$count = 31478;
	#10 counter$count = 31479;
	#10 counter$count = 31480;
	#10 counter$count = 31481;
	#10 counter$count = 31482;
	#10 counter$count = 31483;
	#10 counter$count = 31484;
	#10 counter$count = 31485;
	#10 counter$count = 31486;
	#10 counter$count = 31487;
	#10 counter$count = 31488;
	#10 counter$count = 31489;
	#10 counter$count = 31490;
	#10 counter$count = 31491;
	#10 counter$count = 31492;
	#10 counter$count = 31493;
	#10 counter$count = 31494;
	#10 counter$count = 31495;
	#10 counter$count = 31496;
	#10 counter$count = 31497;
	#10 counter$count = 31498;
	#10 counter$count = 31499;
	#10 counter$count = 31500;
	#10 counter$count = 31501;
	#10 counter$count = 31502;
	#10 counter$count = 31503;
	#10 counter$count = 31504;
	#10 counter$count = 31505;
	#10 counter$count = 31506;
	#10 counter$count = 31507;
	#10 counter$count = 31508;
	#10 counter$count = 31509;
	#10 counter$count = 31510;
	#10 counter$count = 31511;
	#10 counter$count = 31512;
	#10 counter$count = 31513;
	#10 counter$count = 31514;
	#10 counter$count = 31515;
	#10 counter$count = 31516;
	#10 counter$count = 31517;
	#10 counter$count = 31518;
	#10 counter$count = 31519;
	#10 counter$count = 31520;
	#10 counter$count = 31521;
	#10 counter$count = 31522;
	#10 counter$count = 31523;
	#10 counter$count = 31524;
	#10 counter$count = 31525;
	#10 counter$count = 31526;
	#10 counter$count = 31527;
	#10 counter$count = 31528;
	#10 counter$count = 31529;
	#10 counter$count = 31530;
	#10 counter$count = 31531;
	#10 counter$count = 31532;
	#10 counter$count = 31533;
	#10 counter$count = 31534;
	#10 counter$count = 31535;
	#10 counter$count = 31536;
	#10 counter$count = 31537;
	#10 counter$count = 31538;
	#10 counter$count = 31539;
	#10 counter$count = 31540;
	#10 counter$count = 31541;
	#10 counter$count = 31542;
	#10 counter$count = 31543;
	#10 counter$count = 31544;
	#10 counter$count = 31545;
	#10 counter$count = 31546;
	#10 counter$count = 31547;
	#10 counter$count = 31548;
	#10 counter$count = 31549;
	#10 counter$count = 31550;
	#10 counter$count = 31551;
	#10 counter$count = 31552;
	#10 counter$count = 31553;
	#10 counter$count = 31554;
	#10 counter$count = 31555;
	#10 counter$count = 31556;
	#10 counter$count = 31557;
	#10 counter$count = 31558;
	#10 counter$count = 31559;
	#10 counter$count = 31560;
	#10 counter$count = 31561;
	#10 counter$count = 31562;
	#10 counter$count = 31563;
	#10 counter$count = 31564;
	#10 counter$count = 31565;
	#10 counter$count = 31566;
	#10 counter$count = 31567;
	#10 counter$count = 31568;
	#10 counter$count = 31569;
	#10 counter$count = 31570;
	#10 counter$count = 31571;
	#10 counter$count = 31572;
	#10 counter$count = 31573;
	#10 counter$count = 31574;
	#10 counter$count = 31575;
	#10 counter$count = 31576;
	#10 counter$count = 31577;
	#10 counter$count = 31578;
	#10 counter$count = 31579;
	#10 counter$count = 31580;
	#10 counter$count = 31581;
	#10 counter$count = 31582;
	#10 counter$count = 31583;
	#10 counter$count = 31584;
	#10 counter$count = 31585;
	#10 counter$count = 31586;
	#10 counter$count = 31587;
	#10 counter$count = 31588;
	#10 counter$count = 31589;
	#10 counter$count = 31590;
	#10 counter$count = 31591;
	#10 counter$count = 31592;
	#10 counter$count = 31593;
	#10 counter$count = 31594;
	#10 counter$count = 31595;
	#10 counter$count = 31596;
	#10 counter$count = 31597;
	#10 counter$count = 31598;
	#10 counter$count = 31599;
	#10 counter$count = 31600;
	#10 counter$count = 31601;
	#10 counter$count = 31602;
	#10 counter$count = 31603;
	#10 counter$count = 31604;
	#10 counter$count = 31605;
	#10 counter$count = 31606;
	#10 counter$count = 31607;
	#10 counter$count = 31608;
	#10 counter$count = 31609;
	#10 counter$count = 31610;
	#10 counter$count = 31611;
	#10 counter$count = 31612;
	#10 counter$count = 31613;
	#10 counter$count = 31614;
	#10 counter$count = 31615;
	#10 counter$count = 31616;
	#10 counter$count = 31617;
	#10 counter$count = 31618;
	#10 counter$count = 31619;
	#10 counter$count = 31620;
	#10 counter$count = 31621;
	#10 counter$count = 31622;
	#10 counter$count = 31623;
	#10 counter$count = 31624;
	#10 counter$count = 31625;
	#10 counter$count = 31626;
	#10 counter$count = 31627;
	#10 counter$count = 31628;
	#10 counter$count = 31629;
	#10 counter$count = 31630;
	#10 counter$count = 31631;
	#10 counter$count = 31632;
	#10 counter$count = 31633;
	#10 counter$count = 31634;
	#10 counter$count = 31635;
	#10 counter$count = 31636;
	#10 counter$count = 31637;
	#10 counter$count = 31638;
	#10 counter$count = 31639;
	#10 counter$count = 31640;
	#10 counter$count = 31641;
	#10 counter$count = 31642;
	#10 counter$count = 31643;
	#10 counter$count = 31644;
	#10 counter$count = 31645;
	#10 counter$count = 31646;
	#10 counter$count = 31647;
	#10 counter$count = 31648;
	#10 counter$count = 31649;
	#10 counter$count = 31650;
	#10 counter$count = 31651;
	#10 counter$count = 31652;
	#10 counter$count = 31653;
	#10 counter$count = 31654;
	#10 counter$count = 31655;
	#10 counter$count = 31656;
	#10 counter$count = 31657;
	#10 counter$count = 31658;
	#10 counter$count = 31659;
	#10 counter$count = 31660;
	#10 counter$count = 31661;
	#10 counter$count = 31662;
	#10 counter$count = 31663;
	#10 counter$count = 31664;
	#10 counter$count = 31665;
	#10 counter$count = 31666;
	#10 counter$count = 31667;
	#10 counter$count = 31668;
	#10 counter$count = 31669;
	#10 counter$count = 31670;
	#10 counter$count = 31671;
	#10 counter$count = 31672;
	#10 counter$count = 31673;
	#10 counter$count = 31674;
	#10 counter$count = 31675;
	#10 counter$count = 31676;
	#10 counter$count = 31677;
	#10 counter$count = 31678;
	#10 counter$count = 31679;
	#10 counter$count = 31680;
	#10 counter$count = 31681;
	#10 counter$count = 31682;
	#10 counter$count = 31683;
	#10 counter$count = 31684;
	#10 counter$count = 31685;
	#10 counter$count = 31686;
	#10 counter$count = 31687;
	#10 counter$count = 31688;
	#10 counter$count = 31689;
	#10 counter$count = 31690;
	#10 counter$count = 31691;
	#10 counter$count = 31692;
	#10 counter$count = 31693;
	#10 counter$count = 31694;
	#10 counter$count = 31695;
	#10 counter$count = 31696;
	#10 counter$count = 31697;
	#10 counter$count = 31698;
	#10 counter$count = 31699;
	#10 counter$count = 31700;
	#10 counter$count = 31701;
	#10 counter$count = 31702;
	#10 counter$count = 31703;
	#10 counter$count = 31704;
	#10 counter$count = 31705;
	#10 counter$count = 31706;
	#10 counter$count = 31707;
	#10 counter$count = 31708;
	#10 counter$count = 31709;
	#10 counter$count = 31710;
	#10 counter$count = 31711;
	#10 counter$count = 31712;
	#10 counter$count = 31713;
	#10 counter$count = 31714;
	#10 counter$count = 31715;
	#10 counter$count = 31716;
	#10 counter$count = 31717;
	#10 counter$count = 31718;
	#10 counter$count = 31719;
	#10 counter$count = 31720;
	#10 counter$count = 31721;
	#10 counter$count = 31722;
	#10 counter$count = 31723;
	#10 counter$count = 31724;
	#10 counter$count = 31725;
	#10 counter$count = 31726;
	#10 counter$count = 31727;
	#10 counter$count = 31728;
	#10 counter$count = 31729;
	#10 counter$count = 31730;
	#10 counter$count = 31731;
	#10 counter$count = 31732;
	#10 counter$count = 31733;
	#10 counter$count = 31734;
	#10 counter$count = 31735;
	#10 counter$count = 31736;
	#10 counter$count = 31737;
	#10 counter$count = 31738;
	#10 counter$count = 31739;
	#10 counter$count = 31740;
	#10 counter$count = 31741;
	#10 counter$count = 31742;
	#10 counter$count = 31743;
	#10 counter$count = 31744;
	#10 counter$count = 31745;
	#10 counter$count = 31746;
	#10 counter$count = 31747;
	#10 counter$count = 31748;
	#10 counter$count = 31749;
	#10 counter$count = 31750;
	#10 counter$count = 31751;
	#10 counter$count = 31752;
	#10 counter$count = 31753;
	#10 counter$count = 31754;
	#10 counter$count = 31755;
	#10 counter$count = 31756;
	#10 counter$count = 31757;
	#10 counter$count = 31758;
	#10 counter$count = 31759;
	#10 counter$count = 31760;
	#10 counter$count = 31761;
	#10 counter$count = 31762;
	#10 counter$count = 31763;
	#10 counter$count = 31764;
	#10 counter$count = 31765;
	#10 counter$count = 31766;
	#10 counter$count = 31767;
	#10 counter$count = 31768;
	#10 counter$count = 31769;
	#10 counter$count = 31770;
	#10 counter$count = 31771;
	#10 counter$count = 31772;
	#10 counter$count = 31773;
	#10 counter$count = 31774;
	#10 counter$count = 31775;
	#10 counter$count = 31776;
	#10 counter$count = 31777;
	#10 counter$count = 31778;
	#10 counter$count = 31779;
	#10 counter$count = 31780;
	#10 counter$count = 31781;
	#10 counter$count = 31782;
	#10 counter$count = 31783;
	#10 counter$count = 31784;
	#10 counter$count = 31785;
	#10 counter$count = 31786;
	#10 counter$count = 31787;
	#10 counter$count = 31788;
	#10 counter$count = 31789;
	#10 counter$count = 31790;
	#10 counter$count = 31791;
	#10 counter$count = 31792;
	#10 counter$count = 31793;
	#10 counter$count = 31794;
	#10 counter$count = 31795;
	#10 counter$count = 31796;
	#10 counter$count = 31797;
	#10 counter$count = 31798;
	#10 counter$count = 31799;
	#10 counter$count = 31800;
	#10 counter$count = 31801;
	#10 counter$count = 31802;
	#10 counter$count = 31803;
	#10 counter$count = 31804;
	#10 counter$count = 31805;
	#10 counter$count = 31806;
	#10 counter$count = 31807;
	#10 counter$count = 31808;
	#10 counter$count = 31809;
	#10 counter$count = 31810;
	#10 counter$count = 31811;
	#10 counter$count = 31812;
	#10 counter$count = 31813;
	#10 counter$count = 31814;
	#10 counter$count = 31815;
	#10 counter$count = 31816;
	#10 counter$count = 31817;
	#10 counter$count = 31818;
	#10 counter$count = 31819;
	#10 counter$count = 31820;
	#10 counter$count = 31821;
	#10 counter$count = 31822;
	#10 counter$count = 31823;
	#10 counter$count = 31824;
	#10 counter$count = 31825;
	#10 counter$count = 31826;
	#10 counter$count = 31827;
	#10 counter$count = 31828;
	#10 counter$count = 31829;
	#10 counter$count = 31830;
	#10 counter$count = 31831;
	#10 counter$count = 31832;
	#10 counter$count = 31833;
	#10 counter$count = 31834;
	#10 counter$count = 31835;
	#10 counter$count = 31836;
	#10 counter$count = 31837;
	#10 counter$count = 31838;
	#10 counter$count = 31839;
	#10 counter$count = 31840;
	#10 counter$count = 31841;
	#10 counter$count = 31842;
	#10 counter$count = 31843;
	#10 counter$count = 31844;
	#10 counter$count = 31845;
	#10 counter$count = 31846;
	#10 counter$count = 31847;
	#10 counter$count = 31848;
	#10 counter$count = 31849;
	#10 counter$count = 31850;
	#10 counter$count = 31851;
	#10 counter$count = 31852;
	#10 counter$count = 31853;
	#10 counter$count = 31854;
	#10 counter$count = 31855;
	#10 counter$count = 31856;
	#10 counter$count = 31857;
	#10 counter$count = 31858;
	#10 counter$count = 31859;
	#10 counter$count = 31860;
	#10 counter$count = 31861;
	#10 counter$count = 31862;
	#10 counter$count = 31863;
	#10 counter$count = 31864;
	#10 counter$count = 31865;
	#10 counter$count = 31866;
	#10 counter$count = 31867;
	#10 counter$count = 31868;
	#10 counter$count = 31869;
	#10 counter$count = 31870;
	#10 counter$count = 31871;
	#10 counter$count = 31872;
	#10 counter$count = 31873;
	#10 counter$count = 31874;
	#10 counter$count = 31875;
	#10 counter$count = 31876;
	#10 counter$count = 31877;
	#10 counter$count = 31878;
	#10 counter$count = 31879;
	#10 counter$count = 31880;
	#10 counter$count = 31881;
	#10 counter$count = 31882;
	#10 counter$count = 31883;
	#10 counter$count = 31884;
	#10 counter$count = 31885;
	#10 counter$count = 31886;
	#10 counter$count = 31887;
	#10 counter$count = 31888;
	#10 counter$count = 31889;
	#10 counter$count = 31890;
	#10 counter$count = 31891;
	#10 counter$count = 31892;
	#10 counter$count = 31893;
	#10 counter$count = 31894;
	#10 counter$count = 31895;
	#10 counter$count = 31896;
	#10 counter$count = 31897;
	#10 counter$count = 31898;
	#10 counter$count = 31899;
	#10 counter$count = 31900;
	#10 counter$count = 31901;
	#10 counter$count = 31902;
	#10 counter$count = 31903;
	#10 counter$count = 31904;
	#10 counter$count = 31905;
	#10 counter$count = 31906;
	#10 counter$count = 31907;
	#10 counter$count = 31908;
	#10 counter$count = 31909;
	#10 counter$count = 31910;
	#10 counter$count = 31911;
	#10 counter$count = 31912;
	#10 counter$count = 31913;
	#10 counter$count = 31914;
	#10 counter$count = 31915;
	#10 counter$count = 31916;
	#10 counter$count = 31917;
	#10 counter$count = 31918;
	#10 counter$count = 31919;
	#10 counter$count = 31920;
	#10 counter$count = 31921;
	#10 counter$count = 31922;
	#10 counter$count = 31923;
	#10 counter$count = 31924;
	#10 counter$count = 31925;
	#10 counter$count = 31926;
	#10 counter$count = 31927;
	#10 counter$count = 31928;
	#10 counter$count = 31929;
	#10 counter$count = 31930;
	#10 counter$count = 31931;
	#10 counter$count = 31932;
	#10 counter$count = 31933;
	#10 counter$count = 31934;
	#10 counter$count = 31935;
	#10 counter$count = 31936;
	#10 counter$count = 31937;
	#10 counter$count = 31938;
	#10 counter$count = 31939;
	#10 counter$count = 31940;
	#10 counter$count = 31941;
	#10 counter$count = 31942;
	#10 counter$count = 31943;
	#10 counter$count = 31944;
	#10 counter$count = 31945;
	#10 counter$count = 31946;
	#10 counter$count = 31947;
	#10 counter$count = 31948;
	#10 counter$count = 31949;
	#10 counter$count = 31950;
	#10 counter$count = 31951;
	#10 counter$count = 31952;
	#10 counter$count = 31953;
	#10 counter$count = 31954;
	#10 counter$count = 31955;
	#10 counter$count = 31956;
	#10 counter$count = 31957;
	#10 counter$count = 31958;
	#10 counter$count = 31959;
	#10 counter$count = 31960;
	#10 counter$count = 31961;
	#10 counter$count = 31962;
	#10 counter$count = 31963;
	#10 counter$count = 31964;
	#10 counter$count = 31965;
	#10 counter$count = 31966;
	#10 counter$count = 31967;
	#10 counter$count = 31968;
	#10 counter$count = 31969;
	#10 counter$count = 31970;
	#10 counter$count = 31971;
	#10 counter$count = 31972;
	#10 counter$count = 31973;
	#10 counter$count = 31974;
	#10 counter$count = 31975;
	#10 counter$count = 31976;
	#10 counter$count = 31977;
	#10 counter$count = 31978;
	#10 counter$count = 31979;
	#10 counter$count = 31980;
	#10 counter$count = 31981;
	#10 counter$count = 31982;
	#10 counter$count = 31983;
	#10 counter$count = 31984;
	#10 counter$count = 31985;
	#10 counter$count = 31986;
	#10 counter$count = 31987;
	#10 counter$count = 31988;
	#10 counter$count = 31989;
	#10 counter$count = 31990;
	#10 counter$count = 31991;
	#10 counter$count = 31992;
	#10 counter$count = 31993;
	#10 counter$count = 31994;
	#10 counter$count = 31995;
	#10 counter$count = 31996;
	#10 counter$count = 31997;
	#10 counter$count = 31998;
	#10 counter$count = 31999;
	#10 counter$count = 32000;
	#10 counter$count = 32001;
	#10 counter$count = 32002;
	#10 counter$count = 32003;
	#10 counter$count = 32004;
	#10 counter$count = 32005;
	#10 counter$count = 32006;
	#10 counter$count = 32007;
	#10 counter$count = 32008;
	#10 counter$count = 32009;
	#10 counter$count = 32010;
	#10 counter$count = 32011;
	#10 counter$count = 32012;
	#10 counter$count = 32013;
	#10 counter$count = 32014;
	#10 counter$count = 32015;
	#10 counter$count = 32016;
	#10 counter$count = 32017;
	#10 counter$count = 32018;
	#10 counter$count = 32019;
	#10 counter$count = 32020;
	#10 counter$count = 32021;
	#10 counter$count = 32022;
	#10 counter$count = 32023;
	#10 counter$count = 32024;
	#10 counter$count = 32025;
	#10 counter$count = 32026;
	#10 counter$count = 32027;
	#10 counter$count = 32028;
	#10 counter$count = 32029;
	#10 counter$count = 32030;
	#10 counter$count = 32031;
	#10 counter$count = 32032;
	#10 counter$count = 32033;
	#10 counter$count = 32034;
	#10 counter$count = 32035;
	#10 counter$count = 32036;
	#10 counter$count = 32037;
	#10 counter$count = 32038;
	#10 counter$count = 32039;
	#10 counter$count = 32040;
	#10 counter$count = 32041;
	#10 counter$count = 32042;
	#10 counter$count = 32043;
	#10 counter$count = 32044;
	#10 counter$count = 32045;
	#10 counter$count = 32046;
	#10 counter$count = 32047;
	#10 counter$count = 32048;
	#10 counter$count = 32049;
	#10 counter$count = 32050;
	#10 counter$count = 32051;
	#10 counter$count = 32052;
	#10 counter$count = 32053;
	#10 counter$count = 32054;
	#10 counter$count = 32055;
	#10 counter$count = 32056;
	#10 counter$count = 32057;
	#10 counter$count = 32058;
	#10 counter$count = 32059;
	#10 counter$count = 32060;
	#10 counter$count = 32061;
	#10 counter$count = 32062;
	#10 counter$count = 32063;
	#10 counter$count = 32064;
	#10 counter$count = 32065;
	#10 counter$count = 32066;
	#10 counter$count = 32067;
	#10 counter$count = 32068;
	#10 counter$count = 32069;
	#10 counter$count = 32070;
	#10 counter$count = 32071;
	#10 counter$count = 32072;
	#10 counter$count = 32073;
	#10 counter$count = 32074;
	#10 counter$count = 32075;
	#10 counter$count = 32076;
	#10 counter$count = 32077;
	#10 counter$count = 32078;
	#10 counter$count = 32079;
	#10 counter$count = 32080;
	#10 counter$count = 32081;
	#10 counter$count = 32082;
	#10 counter$count = 32083;
	#10 counter$count = 32084;
	#10 counter$count = 32085;
	#10 counter$count = 32086;
	#10 counter$count = 32087;
	#10 counter$count = 32088;
	#10 counter$count = 32089;
	#10 counter$count = 32090;
	#10 counter$count = 32091;
	#10 counter$count = 32092;
	#10 counter$count = 32093;
	#10 counter$count = 32094;
	#10 counter$count = 32095;
	#10 counter$count = 32096;
	#10 counter$count = 32097;
	#10 counter$count = 32098;
	#10 counter$count = 32099;
	#10 counter$count = 32100;
	#10 counter$count = 32101;
	#10 counter$count = 32102;
	#10 counter$count = 32103;
	#10 counter$count = 32104;
	#10 counter$count = 32105;
	#10 counter$count = 32106;
	#10 counter$count = 32107;
	#10 counter$count = 32108;
	#10 counter$count = 32109;
	#10 counter$count = 32110;
	#10 counter$count = 32111;
	#10 counter$count = 32112;
	#10 counter$count = 32113;
	#10 counter$count = 32114;
	#10 counter$count = 32115;
	#10 counter$count = 32116;
	#10 counter$count = 32117;
	#10 counter$count = 32118;
	#10 counter$count = 32119;
	#10 counter$count = 32120;
	#10 counter$count = 32121;
	#10 counter$count = 32122;
	#10 counter$count = 32123;
	#10 counter$count = 32124;
	#10 counter$count = 32125;
	#10 counter$count = 32126;
	#10 counter$count = 32127;
	#10 counter$count = 32128;
	#10 counter$count = 32129;
	#10 counter$count = 32130;
	#10 counter$count = 32131;
	#10 counter$count = 32132;
	#10 counter$count = 32133;
	#10 counter$count = 32134;
	#10 counter$count = 32135;
	#10 counter$count = 32136;
	#10 counter$count = 32137;
	#10 counter$count = 32138;
	#10 counter$count = 32139;
	#10 counter$count = 32140;
	#10 counter$count = 32141;
	#10 counter$count = 32142;
	#10 counter$count = 32143;
	#10 counter$count = 32144;
	#10 counter$count = 32145;
	#10 counter$count = 32146;
	#10 counter$count = 32147;
	#10 counter$count = 32148;
	#10 counter$count = 32149;
	#10 counter$count = 32150;
	#10 counter$count = 32151;
	#10 counter$count = 32152;
	#10 counter$count = 32153;
	#10 counter$count = 32154;
	#10 counter$count = 32155;
	#10 counter$count = 32156;
	#10 counter$count = 32157;
	#10 counter$count = 32158;
	#10 counter$count = 32159;
	#10 counter$count = 32160;
	#10 counter$count = 32161;
	#10 counter$count = 32162;
	#10 counter$count = 32163;
	#10 counter$count = 32164;
	#10 counter$count = 32165;
	#10 counter$count = 32166;
	#10 counter$count = 32167;
	#10 counter$count = 32168;
	#10 counter$count = 32169;
	#10 counter$count = 32170;
	#10 counter$count = 32171;
	#10 counter$count = 32172;
	#10 counter$count = 32173;
	#10 counter$count = 32174;
	#10 counter$count = 32175;
	#10 counter$count = 32176;
	#10 counter$count = 32177;
	#10 counter$count = 32178;
	#10 counter$count = 32179;
	#10 counter$count = 32180;
	#10 counter$count = 32181;
	#10 counter$count = 32182;
	#10 counter$count = 32183;
	#10 counter$count = 32184;
	#10 counter$count = 32185;
	#10 counter$count = 32186;
	#10 counter$count = 32187;
	#10 counter$count = 32188;
	#10 counter$count = 32189;
	#10 counter$count = 32190;
	#10 counter$count = 32191;
	#10 counter$count = 32192;
	#10 counter$count = 32193;
	#10 counter$count = 32194;
	#10 counter$count = 32195;
	#10 counter$count = 32196;
	#10 counter$count = 32197;
	#10 counter$count = 32198;
	#10 counter$count = 32199;
	#10 counter$count = 32200;
	#10 counter$count = 32201;
	#10 counter$count = 32202;
	#10 counter$count = 32203;
	#10 counter$count = 32204;
	#10 counter$count = 32205;
	#10 counter$count = 32206;
	#10 counter$count = 32207;
	#10 counter$count = 32208;
	#10 counter$count = 32209;
	#10 counter$count = 32210;
	#10 counter$count = 32211;
	#10 counter$count = 32212;
	#10 counter$count = 32213;
	#10 counter$count = 32214;
	#10 counter$count = 32215;
	#10 counter$count = 32216;
	#10 counter$count = 32217;
	#10 counter$count = 32218;
	#10 counter$count = 32219;
	#10 counter$count = 32220;
	#10 counter$count = 32221;
	#10 counter$count = 32222;
	#10 counter$count = 32223;
	#10 counter$count = 32224;
	#10 counter$count = 32225;
	#10 counter$count = 32226;
	#10 counter$count = 32227;
	#10 counter$count = 32228;
	#10 counter$count = 32229;
	#10 counter$count = 32230;
	#10 counter$count = 32231;
	#10 counter$count = 32232;
	#10 counter$count = 32233;
	#10 counter$count = 32234;
	#10 counter$count = 32235;
	#10 counter$count = 32236;
	#10 counter$count = 32237;
	#10 counter$count = 32238;
	#10 counter$count = 32239;
	#10 counter$count = 32240;
	#10 counter$count = 32241;
	#10 counter$count = 32242;
	#10 counter$count = 32243;
	#10 counter$count = 32244;
	#10 counter$count = 32245;
	#10 counter$count = 32246;
	#10 counter$count = 32247;
	#10 counter$count = 32248;
	#10 counter$count = 32249;
	#10 counter$count = 32250;
	#10 counter$count = 32251;
	#10 counter$count = 32252;
	#10 counter$count = 32253;
	#10 counter$count = 32254;
	#10 counter$count = 32255;
	#10 counter$count = 32256;
	#10 counter$count = 32257;
	#10 counter$count = 32258;
	#10 counter$count = 32259;
	#10 counter$count = 32260;
	#10 counter$count = 32261;
	#10 counter$count = 32262;
	#10 counter$count = 32263;
	#10 counter$count = 32264;
	#10 counter$count = 32265;
	#10 counter$count = 32266;
	#10 counter$count = 32267;
	#10 counter$count = 32268;
	#10 counter$count = 32269;
	#10 counter$count = 32270;
	#10 counter$count = 32271;
	#10 counter$count = 32272;
	#10 counter$count = 32273;
	#10 counter$count = 32274;
	#10 counter$count = 32275;
	#10 counter$count = 32276;
	#10 counter$count = 32277;
	#10 counter$count = 32278;
	#10 counter$count = 32279;
	#10 counter$count = 32280;
	#10 counter$count = 32281;
	#10 counter$count = 32282;
	#10 counter$count = 32283;
	#10 counter$count = 32284;
	#10 counter$count = 32285;
	#10 counter$count = 32286;
	#10 counter$count = 32287;
	#10 counter$count = 32288;
	#10 counter$count = 32289;
	#10 counter$count = 32290;
	#10 counter$count = 32291;
	#10 counter$count = 32292;
	#10 counter$count = 32293;
	#10 counter$count = 32294;
	#10 counter$count = 32295;
	#10 counter$count = 32296;
	#10 counter$count = 32297;
	#10 counter$count = 32298;
	#10 counter$count = 32299;
	#10 counter$count = 32300;
	#10 counter$count = 32301;
	#10 counter$count = 32302;
	#10 counter$count = 32303;
	#10 counter$count = 32304;
	#10 counter$count = 32305;
	#10 counter$count = 32306;
	#10 counter$count = 32307;
	#10 counter$count = 32308;
	#10 counter$count = 32309;
	#10 counter$count = 32310;
	#10 counter$count = 32311;
	#10 counter$count = 32312;
	#10 counter$count = 32313;
	#10 counter$count = 32314;
	#10 counter$count = 32315;
	#10 counter$count = 32316;
	#10 counter$count = 32317;
	#10 counter$count = 32318;
	#10 counter$count = 32319;
	#10 counter$count = 32320;
	#10 counter$count = 32321;
	#10 counter$count = 32322;
	#10 counter$count = 32323;
	#10 counter$count = 32324;
	#10 counter$count = 32325;
	#10 counter$count = 32326;
	#10 counter$count = 32327;
	#10 counter$count = 32328;
	#10 counter$count = 32329;
	#10 counter$count = 32330;
	#10 counter$count = 32331;
	#10 counter$count = 32332;
	#10 counter$count = 32333;
	#10 counter$count = 32334;
	#10 counter$count = 32335;
	#10 counter$count = 32336;
	#10 counter$count = 32337;
	#10 counter$count = 32338;
	#10 counter$count = 32339;
	#10 counter$count = 32340;
	#10 counter$count = 32341;
	#10 counter$count = 32342;
	#10 counter$count = 32343;
	#10 counter$count = 32344;
	#10 counter$count = 32345;
	#10 counter$count = 32346;
	#10 counter$count = 32347;
	#10 counter$count = 32348;
	#10 counter$count = 32349;
	#10 counter$count = 32350;
	#10 counter$count = 32351;
	#10 counter$count = 32352;
	#10 counter$count = 32353;
	#10 counter$count = 32354;
	#10 counter$count = 32355;
	#10 counter$count = 32356;
	#10 counter$count = 32357;
	#10 counter$count = 32358;
	#10 counter$count = 32359;
	#10 counter$count = 32360;
	#10 counter$count = 32361;
	#10 counter$count = 32362;
	#10 counter$count = 32363;
	#10 counter$count = 32364;
	#10 counter$count = 32365;
	#10 counter$count = 32366;
	#10 counter$count = 32367;
	#10 counter$count = 32368;
	#10 counter$count = 32369;
	#10 counter$count = 32370;
	#10 counter$count = 32371;
	#10 counter$count = 32372;
	#10 counter$count = 32373;
	#10 counter$count = 32374;
	#10 counter$count = 32375;
	#10 counter$count = 32376;
	#10 counter$count = 32377;
	#10 counter$count = 32378;
	#10 counter$count = 32379;
	#10 counter$count = 32380;
	#10 counter$count = 32381;
	#10 counter$count = 32382;
	#10 counter$count = 32383;
	#10 counter$count = 32384;
	#10 counter$count = 32385;
	#10 counter$count = 32386;
	#10 counter$count = 32387;
	#10 counter$count = 32388;
	#10 counter$count = 32389;
	#10 counter$count = 32390;
	#10 counter$count = 32391;
	#10 counter$count = 32392;
	#10 counter$count = 32393;
	#10 counter$count = 32394;
	#10 counter$count = 32395;
	#10 counter$count = 32396;
	#10 counter$count = 32397;
	#10 counter$count = 32398;
	#10 counter$count = 32399;
	#10 counter$count = 32400;
	#10 counter$count = 32401;
	#10 counter$count = 32402;
	#10 counter$count = 32403;
	#10 counter$count = 32404;
	#10 counter$count = 32405;
	#10 counter$count = 32406;
	#10 counter$count = 32407;
	#10 counter$count = 32408;
	#10 counter$count = 32409;
	#10 counter$count = 32410;
	#10 counter$count = 32411;
	#10 counter$count = 32412;
	#10 counter$count = 32413;
	#10 counter$count = 32414;
	#10 counter$count = 32415;
	#10 counter$count = 32416;
	#10 counter$count = 32417;
	#10 counter$count = 32418;
	#10 counter$count = 32419;
	#10 counter$count = 32420;
	#10 counter$count = 32421;
	#10 counter$count = 32422;
	#10 counter$count = 32423;
	#10 counter$count = 32424;
	#10 counter$count = 32425;
	#10 counter$count = 32426;
	#10 counter$count = 32427;
	#10 counter$count = 32428;
	#10 counter$count = 32429;
	#10 counter$count = 32430;
	#10 counter$count = 32431;
	#10 counter$count = 32432;
	#10 counter$count = 32433;
	#10 counter$count = 32434;
	#10 counter$count = 32435;
	#10 counter$count = 32436;
	#10 counter$count = 32437;
	#10 counter$count = 32438;
	#10 counter$count = 32439;
	#10 counter$count = 32440;
	#10 counter$count = 32441;
	#10 counter$count = 32442;
	#10 counter$count = 32443;
	#10 counter$count = 32444;
	#10 counter$count = 32445;
	#10 counter$count = 32446;
	#10 counter$count = 32447;
	#10 counter$count = 32448;
	#10 counter$count = 32449;
	#10 counter$count = 32450;
	#10 counter$count = 32451;
	#10 counter$count = 32452;
	#10 counter$count = 32453;
	#10 counter$count = 32454;
	#10 counter$count = 32455;
	#10 counter$count = 32456;
	#10 counter$count = 32457;
	#10 counter$count = 32458;
	#10 counter$count = 32459;
	#10 counter$count = 32460;
	#10 counter$count = 32461;
	#10 counter$count = 32462;
	#10 counter$count = 32463;
	#10 counter$count = 32464;
	#10 counter$count = 32465;
	#10 counter$count = 32466;
	#10 counter$count = 32467;
	#10 counter$count = 32468;
	#10 counter$count = 32469;
	#10 counter$count = 32470;
	#10 counter$count = 32471;
	#10 counter$count = 32472;
	#10 counter$count = 32473;
	#10 counter$count = 32474;
	#10 counter$count = 32475;
	#10 counter$count = 32476;
	#10 counter$count = 32477;
	#10 counter$count = 32478;
	#10 counter$count = 32479;
	#10 counter$count = 32480;
	#10 counter$count = 32481;
	#10 counter$count = 32482;
	#10 counter$count = 32483;
	#10 counter$count = 32484;
	#10 counter$count = 32485;
	#10 counter$count = 32486;
	#10 counter$count = 32487;
	#10 counter$count = 32488;
	#10 counter$count = 32489;
	#10 counter$count = 32490;
	#10 counter$count = 32491;
	#10 counter$count = 32492;
	#10 counter$count = 32493;
	#10 counter$count = 32494;
	#10 counter$count = 32495;
	#10 counter$count = 32496;
	#10 counter$count = 32497;
	#10 counter$count = 32498;
	#10 counter$count = 32499;
	#10 counter$count = 32500;
	#10 counter$count = 32501;
	#10 counter$count = 32502;
	#10 counter$count = 32503;
	#10 counter$count = 32504;
	#10 counter$count = 32505;
	#10 counter$count = 32506;
	#10 counter$count = 32507;
	#10 counter$count = 32508;
	#10 counter$count = 32509;
	#10 counter$count = 32510;
	#10 counter$count = 32511;
	#10 counter$count = 32512;
	#10 counter$count = 32513;
	#10 counter$count = 32514;
	#10 counter$count = 32515;
	#10 counter$count = 32516;
	#10 counter$count = 32517;
	#10 counter$count = 32518;
	#10 counter$count = 32519;
	#10 counter$count = 32520;
	#10 counter$count = 32521;
	#10 counter$count = 32522;
	#10 counter$count = 32523;
	#10 counter$count = 32524;
	#10 counter$count = 32525;
	#10 counter$count = 32526;
	#10 counter$count = 32527;
	#10 counter$count = 32528;
	#10 counter$count = 32529;
	#10 counter$count = 32530;
	#10 counter$count = 32531;
	#10 counter$count = 32532;
	#10 counter$count = 32533;
	#10 counter$count = 32534;
	#10 counter$count = 32535;
	#10 counter$count = 32536;
	#10 counter$count = 32537;
	#10 counter$count = 32538;
	#10 counter$count = 32539;
	#10 counter$count = 32540;
	#10 counter$count = 32541;
	#10 counter$count = 32542;
	#10 counter$count = 32543;
	#10 counter$count = 32544;
	#10 counter$count = 32545;
	#10 counter$count = 32546;
	#10 counter$count = 32547;
	#10 counter$count = 32548;
	#10 counter$count = 32549;
	#10 counter$count = 32550;
	#10 counter$count = 32551;
	#10 counter$count = 32552;
	#10 counter$count = 32553;
	#10 counter$count = 32554;
	#10 counter$count = 32555;
	#10 counter$count = 32556;
	#10 counter$count = 32557;
	#10 counter$count = 32558;
	#10 counter$count = 32559;
	#10 counter$count = 32560;
	#10 counter$count = 32561;
	#10 counter$count = 32562;
	#10 counter$count = 32563;
	#10 counter$count = 32564;
	#10 counter$count = 32565;
	#10 counter$count = 32566;
	#10 counter$count = 32567;
	#10 counter$count = 32568;
	#10 counter$count = 32569;
	#10 counter$count = 32570;
	#10 counter$count = 32571;
	#10 counter$count = 32572;
	#10 counter$count = 32573;
	#10 counter$count = 32574;
	#10 counter$count = 32575;
	#10 counter$count = 32576;
	#10 counter$count = 32577;
	#10 counter$count = 32578;
	#10 counter$count = 32579;
	#10 counter$count = 32580;
	#10 counter$count = 32581;
	#10 counter$count = 32582;
	#10 counter$count = 32583;
	#10 counter$count = 32584;
	#10 counter$count = 32585;
	#10 counter$count = 32586;
	#10 counter$count = 32587;
	#10 counter$count = 32588;
	#10 counter$count = 32589;
	#10 counter$count = 32590;
	#10 counter$count = 32591;
	#10 counter$count = 32592;
	#10 counter$count = 32593;
	#10 counter$count = 32594;
	#10 counter$count = 32595;
	#10 counter$count = 32596;
	#10 counter$count = 32597;
	#10 counter$count = 32598;
	#10 counter$count = 32599;
	#10 counter$count = 32600;
	#10 counter$count = 32601;
	#10 counter$count = 32602;
	#10 counter$count = 32603;
	#10 counter$count = 32604;
	#10 counter$count = 32605;
	#10 counter$count = 32606;
	#10 counter$count = 32607;
	#10 counter$count = 32608;
	#10 counter$count = 32609;
	#10 counter$count = 32610;
	#10 counter$count = 32611;
	#10 counter$count = 32612;
	#10 counter$count = 32613;
	#10 counter$count = 32614;
	#10 counter$count = 32615;
	#10 counter$count = 32616;
	#10 counter$count = 32617;
	#10 counter$count = 32618;
	#10 counter$count = 32619;
	#10 counter$count = 32620;
	#10 counter$count = 32621;
	#10 counter$count = 32622;
	#10 counter$count = 32623;
	#10 counter$count = 32624;
	#10 counter$count = 32625;
	#10 counter$count = 32626;
	#10 counter$count = 32627;
	#10 counter$count = 32628;
	#10 counter$count = 32629;
	#10 counter$count = 32630;
	#10 counter$count = 32631;
	#10 counter$count = 32632;
	#10 counter$count = 32633;
	#10 counter$count = 32634;
	#10 counter$count = 32635;
	#10 counter$count = 32636;
	#10 counter$count = 32637;
	#10 counter$count = 32638;
	#10 counter$count = 32639;
	#10 counter$count = 32640;
	#10 counter$count = 32641;
	#10 counter$count = 32642;
	#10 counter$count = 32643;
	#10 counter$count = 32644;
	#10 counter$count = 32645;
	#10 counter$count = 32646;
	#10 counter$count = 32647;
	#10 counter$count = 32648;
	#10 counter$count = 32649;
	#10 counter$count = 32650;
	#10 counter$count = 32651;
	#10 counter$count = 32652;
	#10 counter$count = 32653;
	#10 counter$count = 32654;
	#10 counter$count = 32655;
	#10 counter$count = 32656;
	#10 counter$count = 32657;
	#10 counter$count = 32658;
	#10 counter$count = 32659;
	#10 counter$count = 32660;
	#10 counter$count = 32661;
	#10 counter$count = 32662;
	#10 counter$count = 32663;
	#10 counter$count = 32664;
	#10 counter$count = 32665;
	#10 counter$count = 32666;
	#10 counter$count = 32667;
	#10 counter$count = 32668;
	#10 counter$count = 32669;
	#10 counter$count = 32670;
	#10 counter$count = 32671;
	#10 counter$count = 32672;
	#10 counter$count = 32673;
	#10 counter$count = 32674;
	#10 counter$count = 32675;
	#10 counter$count = 32676;
	#10 counter$count = 32677;
	#10 counter$count = 32678;
	#10 counter$count = 32679;
	#10 counter$count = 32680;
	#10 counter$count = 32681;
	#10 counter$count = 32682;
	#10 counter$count = 32683;
	#10 counter$count = 32684;
	#10 counter$count = 32685;
	#10 counter$count = 32686;
	#10 counter$count = 32687;
	#10 counter$count = 32688;
	#10 counter$count = 32689;
	#10 counter$count = 32690;
	#10 counter$count = 32691;
	#10 counter$count = 32692;
	#10 counter$count = 32693;
	#10 counter$count = 32694;
	#10 counter$count = 32695;
	#10 counter$count = 32696;
	#10 counter$count = 32697;
	#10 counter$count = 32698;
	#10 counter$count = 32699;
	#10 counter$count = 32700;
	#10 counter$count = 32701;
	#10 counter$count = 32702;
	#10 counter$count = 32703;
	#10 counter$count = 32704;
	#10 counter$count = 32705;
	#10 counter$count = 32706;
	#10 counter$count = 32707;
	#10 counter$count = 32708;
	#10 counter$count = 32709;
	#10 counter$count = 32710;
	#10 counter$count = 32711;
	#10 counter$count = 32712;
	#10 counter$count = 32713;
	#10 counter$count = 32714;
	#10 counter$count = 32715;
	#10 counter$count = 32716;
	#10 counter$count = 32717;
	#10 counter$count = 32718;
	#10 counter$count = 32719;
	#10 counter$count = 32720;
	#10 counter$count = 32721;
	#10 counter$count = 32722;
	#10 counter$count = 32723;
	#10 counter$count = 32724;
	#10 counter$count = 32725;
	#10 counter$count = 32726;
	#10 counter$count = 32727;
	#10 counter$count = 32728;
	#10 counter$count = 32729;
	#10 counter$count = 32730;
	#10 counter$count = 32731;
	#10 counter$count = 32732;
	#10 counter$count = 32733;
	#10 counter$count = 32734;
	#10 counter$count = 32735;
	#10 counter$count = 32736;
	#10 counter$count = 32737;
	#10 counter$count = 32738;
	#10 counter$count = 32739;
	#10 counter$count = 32740;
	#10 counter$count = 32741;
	#10 counter$count = 32742;
	#10 counter$count = 32743;
	#10 counter$count = 32744;
	#10 counter$count = 32745;
	#10 counter$count = 32746;
	#10 counter$count = 32747;
	#10 counter$count = 32748;
	#10 counter$count = 32749;
	#10 counter$count = 32750;
	#10 counter$count = 32751;
	#10 counter$count = 32752;
	#10 counter$count = 32753;
	#10 counter$count = 32754;
	#10 counter$count = 32755;
	#10 counter$count = 32756;
	#10 counter$count = 32757;
	#10 counter$count = 32758;
	#10 counter$count = 32759;
	#10 counter$count = 32760;
	#10 counter$count = 32761;
	#10 counter$count = 32762;
	#10 counter$count = 32763;
	#10 counter$count = 32764;
	#10 counter$count = 32765;
	#10 counter$count = 32766;
	#10 counter$count = 32767;
	#10 counter$count = 32768;
	#10 counter$count = 32769;
	#10 counter$count = 32770;
	#10 counter$count = 32771;
	#10 counter$count = 32772;
	#10 counter$count = 32773;
	#10 counter$count = 32774;
	#10 counter$count = 32775;
	#10 counter$count = 32776;
	#10 counter$count = 32777;
	#10 counter$count = 32778;
	#10 counter$count = 32779;
	#10 counter$count = 32780;
	#10 counter$count = 32781;
	#10 counter$count = 32782;
	#10 counter$count = 32783;
	#10 counter$count = 32784;
	#10 counter$count = 32785;
	#10 counter$count = 32786;
	#10 counter$count = 32787;
	#10 counter$count = 32788;
	#10 counter$count = 32789;
	#10 counter$count = 32790;
	#10 counter$count = 32791;
	#10 counter$count = 32792;
	#10 counter$count = 32793;
	#10 counter$count = 32794;
	#10 counter$count = 32795;
	#10 counter$count = 32796;
	#10 counter$count = 32797;
	#10 counter$count = 32798;
	#10 counter$count = 32799;
	#10 counter$count = 32800;
	#10 counter$count = 32801;
	#10 counter$count = 32802;
	#10 counter$count = 32803;
	#10 counter$count = 32804;
	#10 counter$count = 32805;
	#10 counter$count = 32806;
	#10 counter$count = 32807;
	#10 counter$count = 32808;
	#10 counter$count = 32809;
	#10 counter$count = 32810;
	#10 counter$count = 32811;
	#10 counter$count = 32812;
	#10 counter$count = 32813;
	#10 counter$count = 32814;
	#10 counter$count = 32815;
	#10 counter$count = 32816;
	#10 counter$count = 32817;
	#10 counter$count = 32818;
	#10 counter$count = 32819;
	#10 counter$count = 32820;
	#10 counter$count = 32821;
	#10 counter$count = 32822;
	#10 counter$count = 32823;
	#10 counter$count = 32824;
	#10 counter$count = 32825;
	#10 counter$count = 32826;
	#10 counter$count = 32827;
	#10 counter$count = 32828;
	#10 counter$count = 32829;
	#10 counter$count = 32830;
	#10 counter$count = 32831;
	#10 counter$count = 32832;
	#10 counter$count = 32833;
	#10 counter$count = 32834;
	#10 counter$count = 32835;
	#10 counter$count = 32836;
	#10 counter$count = 32837;
	#10 counter$count = 32838;
	#10 counter$count = 32839;
	#10 counter$count = 32840;
	#10 counter$count = 32841;
	#10 counter$count = 32842;
	#10 counter$count = 32843;
	#10 counter$count = 32844;
	#10 counter$count = 32845;
	#10 counter$count = 32846;
	#10 counter$count = 32847;
	#10 counter$count = 32848;
	#10 counter$count = 32849;
	#10 counter$count = 32850;
	#10 counter$count = 32851;
	#10 counter$count = 32852;
	#10 counter$count = 32853;
	#10 counter$count = 32854;
	#10 counter$count = 32855;
	#10 counter$count = 32856;
	#10 counter$count = 32857;
	#10 counter$count = 32858;
	#10 counter$count = 32859;
	#10 counter$count = 32860;
	#10 counter$count = 32861;
	#10 counter$count = 32862;
	#10 counter$count = 32863;
	#10 counter$count = 32864;
	#10 counter$count = 32865;
	#10 counter$count = 32866;
	#10 counter$count = 32867;
	#10 counter$count = 32868;
	#10 counter$count = 32869;
	#10 counter$count = 32870;
	#10 counter$count = 32871;
	#10 counter$count = 32872;
	#10 counter$count = 32873;
	#10 counter$count = 32874;
	#10 counter$count = 32875;
	#10 counter$count = 32876;
	#10 counter$count = 32877;
	#10 counter$count = 32878;
	#10 counter$count = 32879;
	#10 counter$count = 32880;
	#10 counter$count = 32881;
	#10 counter$count = 32882;
	#10 counter$count = 32883;
	#10 counter$count = 32884;
	#10 counter$count = 32885;
	#10 counter$count = 32886;
	#10 counter$count = 32887;
	#10 counter$count = 32888;
	#10 counter$count = 32889;
	#10 counter$count = 32890;
	#10 counter$count = 32891;
	#10 counter$count = 32892;
	#10 counter$count = 32893;
	#10 counter$count = 32894;
	#10 counter$count = 32895;
	#10 counter$count = 32896;
	#10 counter$count = 32897;
	#10 counter$count = 32898;
	#10 counter$count = 32899;
	#10 counter$count = 32900;
	#10 counter$count = 32901;
	#10 counter$count = 32902;
	#10 counter$count = 32903;
	#10 counter$count = 32904;
	#10 counter$count = 32905;
	#10 counter$count = 32906;
	#10 counter$count = 32907;
	#10 counter$count = 32908;
	#10 counter$count = 32909;
	#10 counter$count = 32910;
	#10 counter$count = 32911;
	#10 counter$count = 32912;
	#10 counter$count = 32913;
	#10 counter$count = 32914;
	#10 counter$count = 32915;
	#10 counter$count = 32916;
	#10 counter$count = 32917;
	#10 counter$count = 32918;
	#10 counter$count = 32919;
	#10 counter$count = 32920;
	#10 counter$count = 32921;
	#10 counter$count = 32922;
	#10 counter$count = 32923;
	#10 counter$count = 32924;
	#10 counter$count = 32925;
	#10 counter$count = 32926;
	#10 counter$count = 32927;
	#10 counter$count = 32928;
	#10 counter$count = 32929;
	#10 counter$count = 32930;
	#10 counter$count = 32931;
	#10 counter$count = 32932;
	#10 counter$count = 32933;
	#10 counter$count = 32934;
	#10 counter$count = 32935;
	#10 counter$count = 32936;
	#10 counter$count = 32937;
	#10 counter$count = 32938;
	#10 counter$count = 32939;
	#10 counter$count = 32940;
	#10 counter$count = 32941;
	#10 counter$count = 32942;
	#10 counter$count = 32943;
	#10 counter$count = 32944;
	#10 counter$count = 32945;
	#10 counter$count = 32946;
	#10 counter$count = 32947;
	#10 counter$count = 32948;
	#10 counter$count = 32949;
	#10 counter$count = 32950;
	#10 counter$count = 32951;
	#10 counter$count = 32952;
	#10 counter$count = 32953;
	#10 counter$count = 32954;
	#10 counter$count = 32955;
	#10 counter$count = 32956;
	#10 counter$count = 32957;
	#10 counter$count = 32958;
	#10 counter$count = 32959;
	#10 counter$count = 32960;
	#10 counter$count = 32961;
	#10 counter$count = 32962;
	#10 counter$count = 32963;
	#10 counter$count = 32964;
	#10 counter$count = 32965;
	#10 counter$count = 32966;
	#10 counter$count = 32967;
	#10 counter$count = 32968;
	#10 counter$count = 32969;
	#10 counter$count = 32970;
	#10 counter$count = 32971;
	#10 counter$count = 32972;
	#10 counter$count = 32973;
	#10 counter$count = 32974;
	#10 counter$count = 32975;
	#10 counter$count = 32976;
	#10 counter$count = 32977;
	#10 counter$count = 32978;
	#10 counter$count = 32979;
	#10 counter$count = 32980;
	#10 counter$count = 32981;
	#10 counter$count = 32982;
	#10 counter$count = 32983;
	#10 counter$count = 32984;
	#10 counter$count = 32985;
	#10 counter$count = 32986;
	#10 counter$count = 32987;
	#10 counter$count = 32988;
	#10 counter$count = 32989;
	#10 counter$count = 32990;
	#10 counter$count = 32991;
	#10 counter$count = 32992;
	#10 counter$count = 32993;
	#10 counter$count = 32994;
	#10 counter$count = 32995;
	#10 counter$count = 32996;
	#10 counter$count = 32997;
	#10 counter$count = 32998;
	#10 counter$count = 32999;
	#10 counter$count = 33000;
	#10 counter$count = 33001;
	#10 counter$count = 33002;
	#10 counter$count = 33003;
	#10 counter$count = 33004;
	#10 counter$count = 33005;
	#10 counter$count = 33006;
	#10 counter$count = 33007;
	#10 counter$count = 33008;
	#10 counter$count = 33009;
	#10 counter$count = 33010;
	#10 counter$count = 33011;
	#10 counter$count = 33012;
	#10 counter$count = 33013;
	#10 counter$count = 33014;
	#10 counter$count = 33015;
	#10 counter$count = 33016;
	#10 counter$count = 33017;
	#10 counter$count = 33018;
	#10 counter$count = 33019;
	#10 counter$count = 33020;
	#10 counter$count = 33021;
	#10 counter$count = 33022;
	#10 counter$count = 33023;
	#10 counter$count = 33024;
	#10 counter$count = 33025;
	#10 counter$count = 33026;
	#10 counter$count = 33027;
	#10 counter$count = 33028;
	#10 counter$count = 33029;
	#10 counter$count = 33030;
	#10 counter$count = 33031;
	#10 counter$count = 33032;
	#10 counter$count = 33033;
	#10 counter$count = 33034;
	#10 counter$count = 33035;
	#10 counter$count = 33036;
	#10 counter$count = 33037;
	#10 counter$count = 33038;
	#10 counter$count = 33039;
	#10 counter$count = 33040;
	#10 counter$count = 33041;
	#10 counter$count = 33042;
	#10 counter$count = 33043;
	#10 counter$count = 33044;
	#10 counter$count = 33045;
	#10 counter$count = 33046;
	#10 counter$count = 33047;
	#10 counter$count = 33048;
	#10 counter$count = 33049;
	#10 counter$count = 33050;
	#10 counter$count = 33051;
	#10 counter$count = 33052;
	#10 counter$count = 33053;
	#10 counter$count = 33054;
	#10 counter$count = 33055;
	#10 counter$count = 33056;
	#10 counter$count = 33057;
	#10 counter$count = 33058;
	#10 counter$count = 33059;
	#10 counter$count = 33060;
	#10 counter$count = 33061;
	#10 counter$count = 33062;
	#10 counter$count = 33063;
	#10 counter$count = 33064;
	#10 counter$count = 33065;
	#10 counter$count = 33066;
	#10 counter$count = 33067;
	#10 counter$count = 33068;
	#10 counter$count = 33069;
	#10 counter$count = 33070;
	#10 counter$count = 33071;
	#10 counter$count = 33072;
	#10 counter$count = 33073;
	#10 counter$count = 33074;
	#10 counter$count = 33075;
	#10 counter$count = 33076;
	#10 counter$count = 33077;
	#10 counter$count = 33078;
	#10 counter$count = 33079;
	#10 counter$count = 33080;
	#10 counter$count = 33081;
	#10 counter$count = 33082;
	#10 counter$count = 33083;
	#10 counter$count = 33084;
	#10 counter$count = 33085;
	#10 counter$count = 33086;
	#10 counter$count = 33087;
	#10 counter$count = 33088;
	#10 counter$count = 33089;
	#10 counter$count = 33090;
	#10 counter$count = 33091;
	#10 counter$count = 33092;
	#10 counter$count = 33093;
	#10 counter$count = 33094;
	#10 counter$count = 33095;
	#10 counter$count = 33096;
	#10 counter$count = 33097;
	#10 counter$count = 33098;
	#10 counter$count = 33099;
	#10 counter$count = 33100;
	#10 counter$count = 33101;
	#10 counter$count = 33102;
	#10 counter$count = 33103;
	#10 counter$count = 33104;
	#10 counter$count = 33105;
	#10 counter$count = 33106;
	#10 counter$count = 33107;
	#10 counter$count = 33108;
	#10 counter$count = 33109;
	#10 counter$count = 33110;
	#10 counter$count = 33111;
	#10 counter$count = 33112;
	#10 counter$count = 33113;
	#10 counter$count = 33114;
	#10 counter$count = 33115;
	#10 counter$count = 33116;
	#10 counter$count = 33117;
	#10 counter$count = 33118;
	#10 counter$count = 33119;
	#10 counter$count = 33120;
	#10 counter$count = 33121;
	#10 counter$count = 33122;
	#10 counter$count = 33123;
	#10 counter$count = 33124;
	#10 counter$count = 33125;
	#10 counter$count = 33126;
	#10 counter$count = 33127;
	#10 counter$count = 33128;
	#10 counter$count = 33129;
	#10 counter$count = 33130;
	#10 counter$count = 33131;
	#10 counter$count = 33132;
	#10 counter$count = 33133;
	#10 counter$count = 33134;
	#10 counter$count = 33135;
	#10 counter$count = 33136;
	#10 counter$count = 33137;
	#10 counter$count = 33138;
	#10 counter$count = 33139;
	#10 counter$count = 33140;
	#10 counter$count = 33141;
	#10 counter$count = 33142;
	#10 counter$count = 33143;
	#10 counter$count = 33144;
	#10 counter$count = 33145;
	#10 counter$count = 33146;
	#10 counter$count = 33147;
	#10 counter$count = 33148;
	#10 counter$count = 33149;
	#10 counter$count = 33150;
	#10 counter$count = 33151;
	#10 counter$count = 33152;
	#10 counter$count = 33153;
	#10 counter$count = 33154;
	#10 counter$count = 33155;
	#10 counter$count = 33156;
	#10 counter$count = 33157;
	#10 counter$count = 33158;
	#10 counter$count = 33159;
	#10 counter$count = 33160;
	#10 counter$count = 33161;
	#10 counter$count = 33162;
	#10 counter$count = 33163;
	#10 counter$count = 33164;
	#10 counter$count = 33165;
	#10 counter$count = 33166;
	#10 counter$count = 33167;
	#10 counter$count = 33168;
	#10 counter$count = 33169;
	#10 counter$count = 33170;
	#10 counter$count = 33171;
	#10 counter$count = 33172;
	#10 counter$count = 33173;
	#10 counter$count = 33174;
	#10 counter$count = 33175;
	#10 counter$count = 33176;
	#10 counter$count = 33177;
	#10 counter$count = 33178;
	#10 counter$count = 33179;
	#10 counter$count = 33180;
	#10 counter$count = 33181;
	#10 counter$count = 33182;
	#10 counter$count = 33183;
	#10 counter$count = 33184;
	#10 counter$count = 33185;
	#10 counter$count = 33186;
	#10 counter$count = 33187;
	#10 counter$count = 33188;
	#10 counter$count = 33189;
	#10 counter$count = 33190;
	#10 counter$count = 33191;
	#10 counter$count = 33192;
	#10 counter$count = 33193;
	#10 counter$count = 33194;
	#10 counter$count = 33195;
	#10 counter$count = 33196;
	#10 counter$count = 33197;
	#10 counter$count = 33198;
	#10 counter$count = 33199;
	#10 counter$count = 33200;
	#10 counter$count = 33201;
	#10 counter$count = 33202;
	#10 counter$count = 33203;
	#10 counter$count = 33204;
	#10 counter$count = 33205;
	#10 counter$count = 33206;
	#10 counter$count = 33207;
	#10 counter$count = 33208;
	#10 counter$count = 33209;
	#10 counter$count = 33210;
	#10 counter$count = 33211;
	#10 counter$count = 33212;
	#10 counter$count = 33213;
	#10 counter$count = 33214;
	#10 counter$count = 33215;
	#10 counter$count = 33216;
	#10 counter$count = 33217;
	#10 counter$count = 33218;
	#10 counter$count = 33219;
	#10 counter$count = 33220;
	#10 counter$count = 33221;
	#10 counter$count = 33222;
	#10 counter$count = 33223;
	#10 counter$count = 33224;
	#10 counter$count = 33225;
	#10 counter$count = 33226;
	#10 counter$count = 33227;
	#10 counter$count = 33228;
	#10 counter$count = 33229;
	#10 counter$count = 33230;
	#10 counter$count = 33231;
	#10 counter$count = 33232;
	#10 counter$count = 33233;
	#10 counter$count = 33234;
	#10 counter$count = 33235;
	#10 counter$count = 33236;
	#10 counter$count = 33237;
	#10 counter$count = 33238;
	#10 counter$count = 33239;
	#10 counter$count = 33240;
	#10 counter$count = 33241;
	#10 counter$count = 33242;
	#10 counter$count = 33243;
	#10 counter$count = 33244;
	#10 counter$count = 33245;
	#10 counter$count = 33246;
	#10 counter$count = 33247;
	#10 counter$count = 33248;
	#10 counter$count = 33249;
	#10 counter$count = 33250;
	#10 counter$count = 33251;
	#10 counter$count = 33252;
	#10 counter$count = 33253;
	#10 counter$count = 33254;
	#10 counter$count = 33255;
	#10 counter$count = 33256;
	#10 counter$count = 33257;
	#10 counter$count = 33258;
	#10 counter$count = 33259;
	#10 counter$count = 33260;
	#10 counter$count = 33261;
	#10 counter$count = 33262;
	#10 counter$count = 33263;
	#10 counter$count = 33264;
	#10 counter$count = 33265;
	#10 counter$count = 33266;
	#10 counter$count = 33267;
	#10 counter$count = 33268;
	#10 counter$count = 33269;
	#10 counter$count = 33270;
	#10 counter$count = 33271;
	#10 counter$count = 33272;
	#10 counter$count = 33273;
	#10 counter$count = 33274;
	#10 counter$count = 33275;
	#10 counter$count = 33276;
	#10 counter$count = 33277;
	#10 counter$count = 33278;
	#10 counter$count = 33279;
	#10 counter$count = 33280;
	#10 counter$count = 33281;
	#10 counter$count = 33282;
	#10 counter$count = 33283;
	#10 counter$count = 33284;
	#10 counter$count = 33285;
	#10 counter$count = 33286;
	#10 counter$count = 33287;
	#10 counter$count = 33288;
	#10 counter$count = 33289;
	#10 counter$count = 33290;
	#10 counter$count = 33291;
	#10 counter$count = 33292;
	#10 counter$count = 33293;
	#10 counter$count = 33294;
	#10 counter$count = 33295;
	#10 counter$count = 33296;
	#10 counter$count = 33297;
	#10 counter$count = 33298;
	#10 counter$count = 33299;
	#10 counter$count = 33300;
	#10 counter$count = 33301;
	#10 counter$count = 33302;
	#10 counter$count = 33303;
	#10 counter$count = 33304;
	#10 counter$count = 33305;
	#10 counter$count = 33306;
	#10 counter$count = 33307;
	#10 counter$count = 33308;
	#10 counter$count = 33309;
	#10 counter$count = 33310;
	#10 counter$count = 33311;
	#10 counter$count = 33312;
	#10 counter$count = 33313;
	#10 counter$count = 33314;
	#10 counter$count = 33315;
	#10 counter$count = 33316;
	#10 counter$count = 33317;
	#10 counter$count = 33318;
	#10 counter$count = 33319;
	#10 counter$count = 33320;
	#10 counter$count = 33321;
	#10 counter$count = 33322;
	#10 counter$count = 33323;
	#10 counter$count = 33324;
	#10 counter$count = 33325;
	#10 counter$count = 33326;
	#10 counter$count = 33327;
	#10 counter$count = 33328;
	#10 counter$count = 33329;
	#10 counter$count = 33330;
	#10 counter$count = 33331;
	#10 counter$count = 33332;
	#10 counter$count = 33333;
	#10 counter$count = 33334;
	#10 counter$count = 33335;
	#10 counter$count = 33336;
	#10 counter$count = 33337;
	#10 counter$count = 33338;
	#10 counter$count = 33339;
	#10 counter$count = 33340;
	#10 counter$count = 33341;
	#10 counter$count = 33342;
	#10 counter$count = 33343;
	#10 counter$count = 33344;
	#10 counter$count = 33345;
	#10 counter$count = 33346;
	#10 counter$count = 33347;
	#10 counter$count = 33348;
	#10 counter$count = 33349;
	#10 counter$count = 33350;
	#10 counter$count = 33351;
	#10 counter$count = 33352;
	#10 counter$count = 33353;
	#10 counter$count = 33354;
	#10 counter$count = 33355;
	#10 counter$count = 33356;
	#10 counter$count = 33357;
	#10 counter$count = 33358;
	#10 counter$count = 33359;
	#10 counter$count = 33360;
	#10 counter$count = 33361;
	#10 counter$count = 33362;
	#10 counter$count = 33363;
	#10 counter$count = 33364;
	#10 counter$count = 33365;
	#10 counter$count = 33366;
	#10 counter$count = 33367;
	#10 counter$count = 33368;
	#10 counter$count = 33369;
	#10 counter$count = 33370;
	#10 counter$count = 33371;
	#10 counter$count = 33372;
	#10 counter$count = 33373;
	#10 counter$count = 33374;
	#10 counter$count = 33375;
	#10 counter$count = 33376;
	#10 counter$count = 33377;
	#10 counter$count = 33378;
	#10 counter$count = 33379;
	#10 counter$count = 33380;
	#10 counter$count = 33381;
	#10 counter$count = 33382;
	#10 counter$count = 33383;
	#10 counter$count = 33384;
	#10 counter$count = 33385;
	#10 counter$count = 33386;
	#10 counter$count = 33387;
	#10 counter$count = 33388;
	#10 counter$count = 33389;
	#10 counter$count = 33390;
	#10 counter$count = 33391;
	#10 counter$count = 33392;
	#10 counter$count = 33393;
	#10 counter$count = 33394;
	#10 counter$count = 33395;
	#10 counter$count = 33396;
	#10 counter$count = 33397;
	#10 counter$count = 33398;
	#10 counter$count = 33399;
	#10 counter$count = 33400;
	#10 counter$count = 33401;
	#10 counter$count = 33402;
	#10 counter$count = 33403;
	#10 counter$count = 33404;
	#10 counter$count = 33405;
	#10 counter$count = 33406;
	#10 counter$count = 33407;
	#10 counter$count = 33408;
	#10 counter$count = 33409;
	#10 counter$count = 33410;
	#10 counter$count = 33411;
	#10 counter$count = 33412;
	#10 counter$count = 33413;
	#10 counter$count = 33414;
	#10 counter$count = 33415;
	#10 counter$count = 33416;
	#10 counter$count = 33417;
	#10 counter$count = 33418;
	#10 counter$count = 33419;
	#10 counter$count = 33420;
	#10 counter$count = 33421;
	#10 counter$count = 33422;
	#10 counter$count = 33423;
	#10 counter$count = 33424;
	#10 counter$count = 33425;
	#10 counter$count = 33426;
	#10 counter$count = 33427;
	#10 counter$count = 33428;
	#10 counter$count = 33429;
	#10 counter$count = 33430;
	#10 counter$count = 33431;
	#10 counter$count = 33432;
	#10 counter$count = 33433;
	#10 counter$count = 33434;
	#10 counter$count = 33435;
	#10 counter$count = 33436;
	#10 counter$count = 33437;
	#10 counter$count = 33438;
	#10 counter$count = 33439;
	#10 counter$count = 33440;
	#10 counter$count = 33441;
	#10 counter$count = 33442;
	#10 counter$count = 33443;
	#10 counter$count = 33444;
	#10 counter$count = 33445;
	#10 counter$count = 33446;
	#10 counter$count = 33447;
	#10 counter$count = 33448;
	#10 counter$count = 33449;
	#10 counter$count = 33450;
	#10 counter$count = 33451;
	#10 counter$count = 33452;
	#10 counter$count = 33453;
	#10 counter$count = 33454;
	#10 counter$count = 33455;
	#10 counter$count = 33456;
	#10 counter$count = 33457;
	#10 counter$count = 33458;
	#10 counter$count = 33459;
	#10 counter$count = 33460;
	#10 counter$count = 33461;
	#10 counter$count = 33462;
	#10 counter$count = 33463;
	#10 counter$count = 33464;
	#10 counter$count = 33465;
	#10 counter$count = 33466;
	#10 counter$count = 33467;
	#10 counter$count = 33468;
	#10 counter$count = 33469;
	#10 counter$count = 33470;
	#10 counter$count = 33471;
	#10 counter$count = 33472;
	#10 counter$count = 33473;
	#10 counter$count = 33474;
	#10 counter$count = 33475;
	#10 counter$count = 33476;
	#10 counter$count = 33477;
	#10 counter$count = 33478;
	#10 counter$count = 33479;
	#10 counter$count = 33480;
	#10 counter$count = 33481;
	#10 counter$count = 33482;
	#10 counter$count = 33483;
	#10 counter$count = 33484;
	#10 counter$count = 33485;
	#10 counter$count = 33486;
	#10 counter$count = 33487;
	#10 counter$count = 33488;
	#10 counter$count = 33489;
	#10 counter$count = 33490;
	#10 counter$count = 33491;
	#10 counter$count = 33492;
	#10 counter$count = 33493;
	#10 counter$count = 33494;
	#10 counter$count = 33495;
	#10 counter$count = 33496;
	#10 counter$count = 33497;
	#10 counter$count = 33498;
	#10 counter$count = 33499;
	#10 counter$count = 33500;
	#10 counter$count = 33501;
	#10 counter$count = 33502;
	#10 counter$count = 33503;
	#10 counter$count = 33504;
	#10 counter$count = 33505;
	#10 counter$count = 33506;
	#10 counter$count = 33507;
	#10 counter$count = 33508;
	#10 counter$count = 33509;
	#10 counter$count = 33510;
	#10 counter$count = 33511;
	#10 counter$count = 33512;
	#10 counter$count = 33513;
	#10 counter$count = 33514;
	#10 counter$count = 33515;
	#10 counter$count = 33516;
	#10 counter$count = 33517;
	#10 counter$count = 33518;
	#10 counter$count = 33519;
	#10 counter$count = 33520;
	#10 counter$count = 33521;
	#10 counter$count = 33522;
	#10 counter$count = 33523;
	#10 counter$count = 33524;
	#10 counter$count = 33525;
	#10 counter$count = 33526;
	#10 counter$count = 33527;
	#10 counter$count = 33528;
	#10 counter$count = 33529;
	#10 counter$count = 33530;
	#10 counter$count = 33531;
	#10 counter$count = 33532;
	#10 counter$count = 33533;
	#10 counter$count = 33534;
	#10 counter$count = 33535;
	#10 counter$count = 33536;
	#10 counter$count = 33537;
	#10 counter$count = 33538;
	#10 counter$count = 33539;
	#10 counter$count = 33540;
	#10 counter$count = 33541;
	#10 counter$count = 33542;
	#10 counter$count = 33543;
	#10 counter$count = 33544;
	#10 counter$count = 33545;
	#10 counter$count = 33546;
	#10 counter$count = 33547;
	#10 counter$count = 33548;
	#10 counter$count = 33549;
	#10 counter$count = 33550;
	#10 counter$count = 33551;
	#10 counter$count = 33552;
	#10 counter$count = 33553;
	#10 counter$count = 33554;
	#10 counter$count = 33555;
	#10 counter$count = 33556;
	#10 counter$count = 33557;
	#10 counter$count = 33558;
	#10 counter$count = 33559;
	#10 counter$count = 33560;
	#10 counter$count = 33561;
	#10 counter$count = 33562;
	#10 counter$count = 33563;
	#10 counter$count = 33564;
	#10 counter$count = 33565;
	#10 counter$count = 33566;
	#10 counter$count = 33567;
	#10 counter$count = 33568;
	#10 counter$count = 33569;
	#10 counter$count = 33570;
	#10 counter$count = 33571;
	#10 counter$count = 33572;
	#10 counter$count = 33573;
	#10 counter$count = 33574;
	#10 counter$count = 33575;
	#10 counter$count = 33576;
	#10 counter$count = 33577;
	#10 counter$count = 33578;
	#10 counter$count = 33579;
	#10 counter$count = 33580;
	#10 counter$count = 33581;
	#10 counter$count = 33582;
	#10 counter$count = 33583;
	#10 counter$count = 33584;
	#10 counter$count = 33585;
	#10 counter$count = 33586;
	#10 counter$count = 33587;
	#10 counter$count = 33588;
	#10 counter$count = 33589;
	#10 counter$count = 33590;
	#10 counter$count = 33591;
	#10 counter$count = 33592;
	#10 counter$count = 33593;
	#10 counter$count = 33594;
	#10 counter$count = 33595;
	#10 counter$count = 33596;
	#10 counter$count = 33597;
	#10 counter$count = 33598;
	#10 counter$count = 33599;
	#10 counter$count = 33600;
	#10 counter$count = 33601;
	#10 counter$count = 33602;
	#10 counter$count = 33603;
	#10 counter$count = 33604;
	#10 counter$count = 33605;
	#10 counter$count = 33606;
	#10 counter$count = 33607;
	#10 counter$count = 33608;
	#10 counter$count = 33609;
	#10 counter$count = 33610;
	#10 counter$count = 33611;
	#10 counter$count = 33612;
	#10 counter$count = 33613;
	#10 counter$count = 33614;
	#10 counter$count = 33615;
	#10 counter$count = 33616;
	#10 counter$count = 33617;
	#10 counter$count = 33618;
	#10 counter$count = 33619;
	#10 counter$count = 33620;
	#10 counter$count = 33621;
	#10 counter$count = 33622;
	#10 counter$count = 33623;
	#10 counter$count = 33624;
	#10 counter$count = 33625;
	#10 counter$count = 33626;
	#10 counter$count = 33627;
	#10 counter$count = 33628;
	#10 counter$count = 33629;
	#10 counter$count = 33630;
	#10 counter$count = 33631;
	#10 counter$count = 33632;
	#10 counter$count = 33633;
	#10 counter$count = 33634;
	#10 counter$count = 33635;
	#10 counter$count = 33636;
	#10 counter$count = 33637;
	#10 counter$count = 33638;
	#10 counter$count = 33639;
	#10 counter$count = 33640;
	#10 counter$count = 33641;
	#10 counter$count = 33642;
	#10 counter$count = 33643;
	#10 counter$count = 33644;
	#10 counter$count = 33645;
	#10 counter$count = 33646;
	#10 counter$count = 33647;
	#10 counter$count = 33648;
	#10 counter$count = 33649;
	#10 counter$count = 33650;
	#10 counter$count = 33651;
	#10 counter$count = 33652;
	#10 counter$count = 33653;
	#10 counter$count = 33654;
	#10 counter$count = 33655;
	#10 counter$count = 33656;
	#10 counter$count = 33657;
	#10 counter$count = 33658;
	#10 counter$count = 33659;
	#10 counter$count = 33660;
	#10 counter$count = 33661;
	#10 counter$count = 33662;
	#10 counter$count = 33663;
	#10 counter$count = 33664;
	#10 counter$count = 33665;
	#10 counter$count = 33666;
	#10 counter$count = 33667;
	#10 counter$count = 33668;
	#10 counter$count = 33669;
	#10 counter$count = 33670;
	#10 counter$count = 33671;
	#10 counter$count = 33672;
	#10 counter$count = 33673;
	#10 counter$count = 33674;
	#10 counter$count = 33675;
	#10 counter$count = 33676;
	#10 counter$count = 33677;
	#10 counter$count = 33678;
	#10 counter$count = 33679;
	#10 counter$count = 33680;
	#10 counter$count = 33681;
	#10 counter$count = 33682;
	#10 counter$count = 33683;
	#10 counter$count = 33684;
	#10 counter$count = 33685;
	#10 counter$count = 33686;
	#10 counter$count = 33687;
	#10 counter$count = 33688;
	#10 counter$count = 33689;
	#10 counter$count = 33690;
	#10 counter$count = 33691;
	#10 counter$count = 33692;
	#10 counter$count = 33693;
	#10 counter$count = 33694;
	#10 counter$count = 33695;
	#10 counter$count = 33696;
	#10 counter$count = 33697;
	#10 counter$count = 33698;
	#10 counter$count = 33699;
	#10 counter$count = 33700;
	#10 counter$count = 33701;
	#10 counter$count = 33702;
	#10 counter$count = 33703;
	#10 counter$count = 33704;
	#10 counter$count = 33705;
	#10 counter$count = 33706;
	#10 counter$count = 33707;
	#10 counter$count = 33708;
	#10 counter$count = 33709;
	#10 counter$count = 33710;
	#10 counter$count = 33711;
	#10 counter$count = 33712;
	#10 counter$count = 33713;
	#10 counter$count = 33714;
	#10 counter$count = 33715;
	#10 counter$count = 33716;
	#10 counter$count = 33717;
	#10 counter$count = 33718;
	#10 counter$count = 33719;
	#10 counter$count = 33720;
	#10 counter$count = 33721;
	#10 counter$count = 33722;
	#10 counter$count = 33723;
	#10 counter$count = 33724;
	#10 counter$count = 33725;
	#10 counter$count = 33726;
	#10 counter$count = 33727;
	#10 counter$count = 33728;
	#10 counter$count = 33729;
	#10 counter$count = 33730;
	#10 counter$count = 33731;
	#10 counter$count = 33732;
	#10 counter$count = 33733;
	#10 counter$count = 33734;
	#10 counter$count = 33735;
	#10 counter$count = 33736;
	#10 counter$count = 33737;
	#10 counter$count = 33738;
	#10 counter$count = 33739;
	#10 counter$count = 33740;
	#10 counter$count = 33741;
	#10 counter$count = 33742;
	#10 counter$count = 33743;
	#10 counter$count = 33744;
	#10 counter$count = 33745;
	#10 counter$count = 33746;
	#10 counter$count = 33747;
	#10 counter$count = 33748;
	#10 counter$count = 33749;
	#10 counter$count = 33750;
	#10 counter$count = 33751;
	#10 counter$count = 33752;
	#10 counter$count = 33753;
	#10 counter$count = 33754;
	#10 counter$count = 33755;
	#10 counter$count = 33756;
	#10 counter$count = 33757;
	#10 counter$count = 33758;
	#10 counter$count = 33759;
	#10 counter$count = 33760;
	#10 counter$count = 33761;
	#10 counter$count = 33762;
	#10 counter$count = 33763;
	#10 counter$count = 33764;
	#10 counter$count = 33765;
	#10 counter$count = 33766;
	#10 counter$count = 33767;
	#10 counter$count = 33768;
	#10 counter$count = 33769;
	#10 counter$count = 33770;
	#10 counter$count = 33771;
	#10 counter$count = 33772;
	#10 counter$count = 33773;
	#10 counter$count = 33774;
	#10 counter$count = 33775;
	#10 counter$count = 33776;
	#10 counter$count = 33777;
	#10 counter$count = 33778;
	#10 counter$count = 33779;
	#10 counter$count = 33780;
	#10 counter$count = 33781;
	#10 counter$count = 33782;
	#10 counter$count = 33783;
	#10 counter$count = 33784;
	#10 counter$count = 33785;
	#10 counter$count = 33786;
	#10 counter$count = 33787;
	#10 counter$count = 33788;
	#10 counter$count = 33789;
	#10 counter$count = 33790;
	#10 counter$count = 33791;
	#10 counter$count = 33792;
	#10 counter$count = 33793;
	#10 counter$count = 33794;
	#10 counter$count = 33795;
	#10 counter$count = 33796;
	#10 counter$count = 33797;
	#10 counter$count = 33798;
	#10 counter$count = 33799;
	#10 counter$count = 33800;
	#10 counter$count = 33801;
	#10 counter$count = 33802;
	#10 counter$count = 33803;
	#10 counter$count = 33804;
	#10 counter$count = 33805;
	#10 counter$count = 33806;
	#10 counter$count = 33807;
	#10 counter$count = 33808;
	#10 counter$count = 33809;
	#10 counter$count = 33810;
	#10 counter$count = 33811;
	#10 counter$count = 33812;
	#10 counter$count = 33813;
	#10 counter$count = 33814;
	#10 counter$count = 33815;
	#10 counter$count = 33816;
	#10 counter$count = 33817;
	#10 counter$count = 33818;
	#10 counter$count = 33819;
	#10 counter$count = 33820;
	#10 counter$count = 33821;
	#10 counter$count = 33822;
	#10 counter$count = 33823;
	#10 counter$count = 33824;
	#10 counter$count = 33825;
	#10 counter$count = 33826;
	#10 counter$count = 33827;
	#10 counter$count = 33828;
	#10 counter$count = 33829;
	#10 counter$count = 33830;
	#10 counter$count = 33831;
	#10 counter$count = 33832;
	#10 counter$count = 33833;
	#10 counter$count = 33834;
	#10 counter$count = 33835;
	#10 counter$count = 33836;
	#10 counter$count = 33837;
	#10 counter$count = 33838;
	#10 counter$count = 33839;
	#10 counter$count = 33840;
	#10 counter$count = 33841;
	#10 counter$count = 33842;
	#10 counter$count = 33843;
	#10 counter$count = 33844;
	#10 counter$count = 33845;
	#10 counter$count = 33846;
	#10 counter$count = 33847;
	#10 counter$count = 33848;
	#10 counter$count = 33849;
	#10 counter$count = 33850;
	#10 counter$count = 33851;
	#10 counter$count = 33852;
	#10 counter$count = 33853;
	#10 counter$count = 33854;
	#10 counter$count = 33855;
	#10 counter$count = 33856;
	#10 counter$count = 33857;
	#10 counter$count = 33858;
	#10 counter$count = 33859;
	#10 counter$count = 33860;
	#10 counter$count = 33861;
	#10 counter$count = 33862;
	#10 counter$count = 33863;
	#10 counter$count = 33864;
	#10 counter$count = 33865;
	#10 counter$count = 33866;
	#10 counter$count = 33867;
	#10 counter$count = 33868;
	#10 counter$count = 33869;
	#10 counter$count = 33870;
	#10 counter$count = 33871;
	#10 counter$count = 33872;
	#10 counter$count = 33873;
	#10 counter$count = 33874;
	#10 counter$count = 33875;
	#10 counter$count = 33876;
	#10 counter$count = 33877;
	#10 counter$count = 33878;
	#10 counter$count = 33879;
	#10 counter$count = 33880;
	#10 counter$count = 33881;
	#10 counter$count = 33882;
	#10 counter$count = 33883;
	#10 counter$count = 33884;
	#10 counter$count = 33885;
	#10 counter$count = 33886;
	#10 counter$count = 33887;
	#10 counter$count = 33888;
	#10 counter$count = 33889;
	#10 counter$count = 33890;
	#10 counter$count = 33891;
	#10 counter$count = 33892;
	#10 counter$count = 33893;
	#10 counter$count = 33894;
	#10 counter$count = 33895;
	#10 counter$count = 33896;
	#10 counter$count = 33897;
	#10 counter$count = 33898;
	#10 counter$count = 33899;
	#10 counter$count = 33900;
	#10 counter$count = 33901;
	#10 counter$count = 33902;
	#10 counter$count = 33903;
	#10 counter$count = 33904;
	#10 counter$count = 33905;
	#10 counter$count = 33906;
	#10 counter$count = 33907;
	#10 counter$count = 33908;
	#10 counter$count = 33909;
	#10 counter$count = 33910;
	#10 counter$count = 33911;
	#10 counter$count = 33912;
	#10 counter$count = 33913;
	#10 counter$count = 33914;
	#10 counter$count = 33915;
	#10 counter$count = 33916;
	#10 counter$count = 33917;
	#10 counter$count = 33918;
	#10 counter$count = 33919;
	#10 counter$count = 33920;
	#10 counter$count = 33921;
	#10 counter$count = 33922;
	#10 counter$count = 33923;
	#10 counter$count = 33924;
	#10 counter$count = 33925;
	#10 counter$count = 33926;
	#10 counter$count = 33927;
	#10 counter$count = 33928;
	#10 counter$count = 33929;
	#10 counter$count = 33930;
	#10 counter$count = 33931;
	#10 counter$count = 33932;
	#10 counter$count = 33933;
	#10 counter$count = 33934;
	#10 counter$count = 33935;
	#10 counter$count = 33936;
	#10 counter$count = 33937;
	#10 counter$count = 33938;
	#10 counter$count = 33939;
	#10 counter$count = 33940;
	#10 counter$count = 33941;
	#10 counter$count = 33942;
	#10 counter$count = 33943;
	#10 counter$count = 33944;
	#10 counter$count = 33945;
	#10 counter$count = 33946;
	#10 counter$count = 33947;
	#10 counter$count = 33948;
	#10 counter$count = 33949;
	#10 counter$count = 33950;
	#10 counter$count = 33951;
	#10 counter$count = 33952;
	#10 counter$count = 33953;
	#10 counter$count = 33954;
	#10 counter$count = 33955;
	#10 counter$count = 33956;
	#10 counter$count = 33957;
	#10 counter$count = 33958;
	#10 counter$count = 33959;
	#10 counter$count = 33960;
	#10 counter$count = 33961;
	#10 counter$count = 33962;
	#10 counter$count = 33963;
	#10 counter$count = 33964;
	#10 counter$count = 33965;
	#10 counter$count = 33966;
	#10 counter$count = 33967;
	#10 counter$count = 33968;
	#10 counter$count = 33969;
	#10 counter$count = 33970;
	#10 counter$count = 33971;
	#10 counter$count = 33972;
	#10 counter$count = 33973;
	#10 counter$count = 33974;
	#10 counter$count = 33975;
	#10 counter$count = 33976;
	#10 counter$count = 33977;
	#10 counter$count = 33978;
	#10 counter$count = 33979;
	#10 counter$count = 33980;
	#10 counter$count = 33981;
	#10 counter$count = 33982;
	#10 counter$count = 33983;
	#10 counter$count = 33984;
	#10 counter$count = 33985;
	#10 counter$count = 33986;
	#10 counter$count = 33987;
	#10 counter$count = 33988;
	#10 counter$count = 33989;
	#10 counter$count = 33990;
	#10 counter$count = 33991;
	#10 counter$count = 33992;
	#10 counter$count = 33993;
	#10 counter$count = 33994;
	#10 counter$count = 33995;
	#10 counter$count = 33996;
	#10 counter$count = 33997;
	#10 counter$count = 33998;
	#10 counter$count = 33999;
	#10 counter$count = 34000;
	#10 counter$count = 34001;
	#10 counter$count = 34002;
	#10 counter$count = 34003;
	#10 counter$count = 34004;
	#10 counter$count = 34005;
	#10 counter$count = 34006;
	#10 counter$count = 34007;
	#10 counter$count = 34008;
	#10 counter$count = 34009;
	#10 counter$count = 34010;
	#10 counter$count = 34011;
	#10 counter$count = 34012;
	#10 counter$count = 34013;
	#10 counter$count = 34014;
	#10 counter$count = 34015;
	#10 counter$count = 34016;
	#10 counter$count = 34017;
	#10 counter$count = 34018;
	#10 counter$count = 34019;
	#10 counter$count = 34020;
	#10 counter$count = 34021;
	#10 counter$count = 34022;
	#10 counter$count = 34023;
	#10 counter$count = 34024;
	#10 counter$count = 34025;
	#10 counter$count = 34026;
	#10 counter$count = 34027;
	#10 counter$count = 34028;
	#10 counter$count = 34029;
	#10 counter$count = 34030;
	#10 counter$count = 34031;
	#10 counter$count = 34032;
	#10 counter$count = 34033;
	#10 counter$count = 34034;
	#10 counter$count = 34035;
	#10 counter$count = 34036;
	#10 counter$count = 34037;
	#10 counter$count = 34038;
	#10 counter$count = 34039;
	#10 counter$count = 34040;
	#10 counter$count = 34041;
	#10 counter$count = 34042;
	#10 counter$count = 34043;
	#10 counter$count = 34044;
	#10 counter$count = 34045;
	#10 counter$count = 34046;
	#10 counter$count = 34047;
	#10 counter$count = 34048;
	#10 counter$count = 34049;
	#10 counter$count = 34050;
	#10 counter$count = 34051;
	#10 counter$count = 34052;
	#10 counter$count = 34053;
	#10 counter$count = 34054;
	#10 counter$count = 34055;
	#10 counter$count = 34056;
	#10 counter$count = 34057;
	#10 counter$count = 34058;
	#10 counter$count = 34059;
	#10 counter$count = 34060;
	#10 counter$count = 34061;
	#10 counter$count = 34062;
	#10 counter$count = 34063;
	#10 counter$count = 34064;
	#10 counter$count = 34065;
	#10 counter$count = 34066;
	#10 counter$count = 34067;
	#10 counter$count = 34068;
	#10 counter$count = 34069;
	#10 counter$count = 34070;
	#10 counter$count = 34071;
	#10 counter$count = 34072;
	#10 counter$count = 34073;
	#10 counter$count = 34074;
	#10 counter$count = 34075;
	#10 counter$count = 34076;
	#10 counter$count = 34077;
	#10 counter$count = 34078;
	#10 counter$count = 34079;
	#10 counter$count = 34080;
	#10 counter$count = 34081;
	#10 counter$count = 34082;
	#10 counter$count = 34083;
	#10 counter$count = 34084;
	#10 counter$count = 34085;
	#10 counter$count = 34086;
	#10 counter$count = 34087;
	#10 counter$count = 34088;
	#10 counter$count = 34089;
	#10 counter$count = 34090;
	#10 counter$count = 34091;
	#10 counter$count = 34092;
	#10 counter$count = 34093;
	#10 counter$count = 34094;
	#10 counter$count = 34095;
	#10 counter$count = 34096;
	#10 counter$count = 34097;
	#10 counter$count = 34098;
	#10 counter$count = 34099;
	#10 counter$count = 34100;
	#10 counter$count = 34101;
	#10 counter$count = 34102;
	#10 counter$count = 34103;
	#10 counter$count = 34104;
	#10 counter$count = 34105;
	#10 counter$count = 34106;
	#10 counter$count = 34107;
	#10 counter$count = 34108;
	#10 counter$count = 34109;
	#10 counter$count = 34110;
	#10 counter$count = 34111;
	#10 counter$count = 34112;
	#10 counter$count = 34113;
	#10 counter$count = 34114;
	#10 counter$count = 34115;
	#10 counter$count = 34116;
	#10 counter$count = 34117;
	#10 counter$count = 34118;
	#10 counter$count = 34119;
	#10 counter$count = 34120;
	#10 counter$count = 34121;
	#10 counter$count = 34122;
	#10 counter$count = 34123;
	#10 counter$count = 34124;
	#10 counter$count = 34125;
	#10 counter$count = 34126;
	#10 counter$count = 34127;
	#10 counter$count = 34128;
	#10 counter$count = 34129;
	#10 counter$count = 34130;
	#10 counter$count = 34131;
	#10 counter$count = 34132;
	#10 counter$count = 34133;
	#10 counter$count = 34134;
	#10 counter$count = 34135;
	#10 counter$count = 34136;
	#10 counter$count = 34137;
	#10 counter$count = 34138;
	#10 counter$count = 34139;
	#10 counter$count = 34140;
	#10 counter$count = 34141;
	#10 counter$count = 34142;
	#10 counter$count = 34143;
	#10 counter$count = 34144;
	#10 counter$count = 34145;
	#10 counter$count = 34146;
	#10 counter$count = 34147;
	#10 counter$count = 34148;
	#10 counter$count = 34149;
	#10 counter$count = 34150;
	#10 counter$count = 34151;
	#10 counter$count = 34152;
	#10 counter$count = 34153;
	#10 counter$count = 34154;
	#10 counter$count = 34155;
	#10 counter$count = 34156;
	#10 counter$count = 34157;
	#10 counter$count = 34158;
	#10 counter$count = 34159;
	#10 counter$count = 34160;
	#10 counter$count = 34161;
	#10 counter$count = 34162;
	#10 counter$count = 34163;
	#10 counter$count = 34164;
	#10 counter$count = 34165;
	#10 counter$count = 34166;
	#10 counter$count = 34167;
	#10 counter$count = 34168;
	#10 counter$count = 34169;
	#10 counter$count = 34170;
	#10 counter$count = 34171;
	#10 counter$count = 34172;
	#10 counter$count = 34173;
	#10 counter$count = 34174;
	#10 counter$count = 34175;
	#10 counter$count = 34176;
	#10 counter$count = 34177;
	#10 counter$count = 34178;
	#10 counter$count = 34179;
	#10 counter$count = 34180;
	#10 counter$count = 34181;
	#10 counter$count = 34182;
	#10 counter$count = 34183;
	#10 counter$count = 34184;
	#10 counter$count = 34185;
	#10 counter$count = 34186;
	#10 counter$count = 34187;
	#10 counter$count = 34188;
	#10 counter$count = 34189;
	#10 counter$count = 34190;
	#10 counter$count = 34191;
	#10 counter$count = 34192;
	#10 counter$count = 34193;
	#10 counter$count = 34194;
	#10 counter$count = 34195;
	#10 counter$count = 34196;
	#10 counter$count = 34197;
	#10 counter$count = 34198;
	#10 counter$count = 34199;
	#10 counter$count = 34200;
	#10 counter$count = 34201;
	#10 counter$count = 34202;
	#10 counter$count = 34203;
	#10 counter$count = 34204;
	#10 counter$count = 34205;
	#10 counter$count = 34206;
	#10 counter$count = 34207;
	#10 counter$count = 34208;
	#10 counter$count = 34209;
	#10 counter$count = 34210;
	#10 counter$count = 34211;
	#10 counter$count = 34212;
	#10 counter$count = 34213;
	#10 counter$count = 34214;
	#10 counter$count = 34215;
	#10 counter$count = 34216;
	#10 counter$count = 34217;
	#10 counter$count = 34218;
	#10 counter$count = 34219;
	#10 counter$count = 34220;
	#10 counter$count = 34221;
	#10 counter$count = 34222;
	#10 counter$count = 34223;
	#10 counter$count = 34224;
	#10 counter$count = 34225;
	#10 counter$count = 34226;
	#10 counter$count = 34227;
	#10 counter$count = 34228;
	#10 counter$count = 34229;
	#10 counter$count = 34230;
	#10 counter$count = 34231;
	#10 counter$count = 34232;
	#10 counter$count = 34233;
	#10 counter$count = 34234;
	#10 counter$count = 34235;
	#10 counter$count = 34236;
	#10 counter$count = 34237;
	#10 counter$count = 34238;
	#10 counter$count = 34239;
	#10 counter$count = 34240;
	#10 counter$count = 34241;
	#10 counter$count = 34242;
	#10 counter$count = 34243;
	#10 counter$count = 34244;
	#10 counter$count = 34245;
	#10 counter$count = 34246;
	#10 counter$count = 34247;
	#10 counter$count = 34248;
	#10 counter$count = 34249;
	#10 counter$count = 34250;
	#10 counter$count = 34251;
	#10 counter$count = 34252;
	#10 counter$count = 34253;
	#10 counter$count = 34254;
	#10 counter$count = 34255;
	#10 counter$count = 34256;
	#10 counter$count = 34257;
	#10 counter$count = 34258;
	#10 counter$count = 34259;
	#10 counter$count = 34260;
	#10 counter$count = 34261;
	#10 counter$count = 34262;
	#10 counter$count = 34263;
	#10 counter$count = 34264;
	#10 counter$count = 34265;
	#10 counter$count = 34266;
	#10 counter$count = 34267;
	#10 counter$count = 34268;
	#10 counter$count = 34269;
	#10 counter$count = 34270;
	#10 counter$count = 34271;
	#10 counter$count = 34272;
	#10 counter$count = 34273;
	#10 counter$count = 34274;
	#10 counter$count = 34275;
	#10 counter$count = 34276;
	#10 counter$count = 34277;
	#10 counter$count = 34278;
	#10 counter$count = 34279;
	#10 counter$count = 34280;
	#10 counter$count = 34281;
	#10 counter$count = 34282;
	#10 counter$count = 34283;
	#10 counter$count = 34284;
	#10 counter$count = 34285;
	#10 counter$count = 34286;
	#10 counter$count = 34287;
	#10 counter$count = 34288;
	#10 counter$count = 34289;
	#10 counter$count = 34290;
	#10 counter$count = 34291;
	#10 counter$count = 34292;
	#10 counter$count = 34293;
	#10 counter$count = 34294;
	#10 counter$count = 34295;
	#10 counter$count = 34296;
	#10 counter$count = 34297;
	#10 counter$count = 34298;
	#10 counter$count = 34299;
	#10 counter$count = 34300;
	#10 counter$count = 34301;
	#10 counter$count = 34302;
	#10 counter$count = 34303;
	#10 counter$count = 34304;
	#10 counter$count = 34305;
	#10 counter$count = 34306;
	#10 counter$count = 34307;
	#10 counter$count = 34308;
	#10 counter$count = 34309;
	#10 counter$count = 34310;
	#10 counter$count = 34311;
	#10 counter$count = 34312;
	#10 counter$count = 34313;
	#10 counter$count = 34314;
	#10 counter$count = 34315;
	#10 counter$count = 34316;
	#10 counter$count = 34317;
	#10 counter$count = 34318;
	#10 counter$count = 34319;
	#10 counter$count = 34320;
	#10 counter$count = 34321;
	#10 counter$count = 34322;
	#10 counter$count = 34323;
	#10 counter$count = 34324;
	#10 counter$count = 34325;
	#10 counter$count = 34326;
	#10 counter$count = 34327;
	#10 counter$count = 34328;
	#10 counter$count = 34329;
	#10 counter$count = 34330;
	#10 counter$count = 34331;
	#10 counter$count = 34332;
	#10 counter$count = 34333;
	#10 counter$count = 34334;
	#10 counter$count = 34335;
	#10 counter$count = 34336;
	#10 counter$count = 34337;
	#10 counter$count = 34338;
	#10 counter$count = 34339;
	#10 counter$count = 34340;
	#10 counter$count = 34341;
	#10 counter$count = 34342;
	#10 counter$count = 34343;
	#10 counter$count = 34344;
	#10 counter$count = 34345;
	#10 counter$count = 34346;
	#10 counter$count = 34347;
	#10 counter$count = 34348;
	#10 counter$count = 34349;
	#10 counter$count = 34350;
	#10 counter$count = 34351;
	#10 counter$count = 34352;
	#10 counter$count = 34353;
	#10 counter$count = 34354;
	#10 counter$count = 34355;
	#10 counter$count = 34356;
	#10 counter$count = 34357;
	#10 counter$count = 34358;
	#10 counter$count = 34359;
	#10 counter$count = 34360;
	#10 counter$count = 34361;
	#10 counter$count = 34362;
	#10 counter$count = 34363;
	#10 counter$count = 34364;
	#10 counter$count = 34365;
	#10 counter$count = 34366;
	#10 counter$count = 34367;
	#10 counter$count = 34368;
	#10 counter$count = 34369;
	#10 counter$count = 34370;
	#10 counter$count = 34371;
	#10 counter$count = 34372;
	#10 counter$count = 34373;
	#10 counter$count = 34374;
	#10 counter$count = 34375;
	#10 counter$count = 34376;
	#10 counter$count = 34377;
	#10 counter$count = 34378;
	#10 counter$count = 34379;
	#10 counter$count = 34380;
	#10 counter$count = 34381;
	#10 counter$count = 34382;
	#10 counter$count = 34383;
	#10 counter$count = 34384;
	#10 counter$count = 34385;
	#10 counter$count = 34386;
	#10 counter$count = 34387;
	#10 counter$count = 34388;
	#10 counter$count = 34389;
	#10 counter$count = 34390;
	#10 counter$count = 34391;
	#10 counter$count = 34392;
	#10 counter$count = 34393;
	#10 counter$count = 34394;
	#10 counter$count = 34395;
	#10 counter$count = 34396;
	#10 counter$count = 34397;
	#10 counter$count = 34398;
	#10 counter$count = 34399;
	#10 counter$count = 34400;
	#10 counter$count = 34401;
	#10 counter$count = 34402;
	#10 counter$count = 34403;
	#10 counter$count = 34404;
	#10 counter$count = 34405;
	#10 counter$count = 34406;
	#10 counter$count = 34407;
	#10 counter$count = 34408;
	#10 counter$count = 34409;
	#10 counter$count = 34410;
	#10 counter$count = 34411;
	#10 counter$count = 34412;
	#10 counter$count = 34413;
	#10 counter$count = 34414;
	#10 counter$count = 34415;
	#10 counter$count = 34416;
	#10 counter$count = 34417;
	#10 counter$count = 34418;
	#10 counter$count = 34419;
	#10 counter$count = 34420;
	#10 counter$count = 34421;
	#10 counter$count = 34422;
	#10 counter$count = 34423;
	#10 counter$count = 34424;
	#10 counter$count = 34425;
	#10 counter$count = 34426;
	#10 counter$count = 34427;
	#10 counter$count = 34428;
	#10 counter$count = 34429;
	#10 counter$count = 34430;
	#10 counter$count = 34431;
	#10 counter$count = 34432;
	#10 counter$count = 34433;
	#10 counter$count = 34434;
	#10 counter$count = 34435;
	#10 counter$count = 34436;
	#10 counter$count = 34437;
	#10 counter$count = 34438;
	#10 counter$count = 34439;
	#10 counter$count = 34440;
	#10 counter$count = 34441;
	#10 counter$count = 34442;
	#10 counter$count = 34443;
	#10 counter$count = 34444;
	#10 counter$count = 34445;
	#10 counter$count = 34446;
	#10 counter$count = 34447;
	#10 counter$count = 34448;
	#10 counter$count = 34449;
	#10 counter$count = 34450;
	#10 counter$count = 34451;
	#10 counter$count = 34452;
	#10 counter$count = 34453;
	#10 counter$count = 34454;
	#10 counter$count = 34455;
	#10 counter$count = 34456;
	#10 counter$count = 34457;
	#10 counter$count = 34458;
	#10 counter$count = 34459;
	#10 counter$count = 34460;
	#10 counter$count = 34461;
	#10 counter$count = 34462;
	#10 counter$count = 34463;
	#10 counter$count = 34464;
	#10 counter$count = 34465;
	#10 counter$count = 34466;
	#10 counter$count = 34467;
	#10 counter$count = 34468;
	#10 counter$count = 34469;
	#10 counter$count = 34470;
	#10 counter$count = 34471;
	#10 counter$count = 34472;
	#10 counter$count = 34473;
	#10 counter$count = 34474;
	#10 counter$count = 34475;
	#10 counter$count = 34476;
	#10 counter$count = 34477;
	#10 counter$count = 34478;
	#10 counter$count = 34479;
	#10 counter$count = 34480;
	#10 counter$count = 34481;
	#10 counter$count = 34482;
	#10 counter$count = 34483;
	#10 counter$count = 34484;
	#10 counter$count = 34485;
	#10 counter$count = 34486;
	#10 counter$count = 34487;
	#10 counter$count = 34488;
	#10 counter$count = 34489;
	#10 counter$count = 34490;
	#10 counter$count = 34491;
	#10 counter$count = 34492;
	#10 counter$count = 34493;
	#10 counter$count = 34494;
	#10 counter$count = 34495;
	#10 counter$count = 34496;
	#10 counter$count = 34497;
	#10 counter$count = 34498;
	#10 counter$count = 34499;
	#10 counter$count = 34500;
	#10 counter$count = 34501;
	#10 counter$count = 34502;
	#10 counter$count = 34503;
	#10 counter$count = 34504;
	#10 counter$count = 34505;
	#10 counter$count = 34506;
	#10 counter$count = 34507;
	#10 counter$count = 34508;
	#10 counter$count = 34509;
	#10 counter$count = 34510;
	#10 counter$count = 34511;
	#10 counter$count = 34512;
	#10 counter$count = 34513;
	#10 counter$count = 34514;
	#10 counter$count = 34515;
	#10 counter$count = 34516;
	#10 counter$count = 34517;
	#10 counter$count = 34518;
	#10 counter$count = 34519;
	#10 counter$count = 34520;
	#10 counter$count = 34521;
	#10 counter$count = 34522;
	#10 counter$count = 34523;
	#10 counter$count = 34524;
	#10 counter$count = 34525;
	#10 counter$count = 34526;
	#10 counter$count = 34527;
	#10 counter$count = 34528;
	#10 counter$count = 34529;
	#10 counter$count = 34530;
	#10 counter$count = 34531;
	#10 counter$count = 34532;
	#10 counter$count = 34533;
	#10 counter$count = 34534;
	#10 counter$count = 34535;
	#10 counter$count = 34536;
	#10 counter$count = 34537;
	#10 counter$count = 34538;
	#10 counter$count = 34539;
	#10 counter$count = 34540;
	#10 counter$count = 34541;
	#10 counter$count = 34542;
	#10 counter$count = 34543;
	#10 counter$count = 34544;
	#10 counter$count = 34545;
	#10 counter$count = 34546;
	#10 counter$count = 34547;
	#10 counter$count = 34548;
	#10 counter$count = 34549;
	#10 counter$count = 34550;
	#10 counter$count = 34551;
	#10 counter$count = 34552;
	#10 counter$count = 34553;
	#10 counter$count = 34554;
	#10 counter$count = 34555;
	#10 counter$count = 34556;
	#10 counter$count = 34557;
	#10 counter$count = 34558;
	#10 counter$count = 34559;
	#10 counter$count = 34560;
	#10 counter$count = 34561;
	#10 counter$count = 34562;
	#10 counter$count = 34563;
	#10 counter$count = 34564;
	#10 counter$count = 34565;
	#10 counter$count = 34566;
	#10 counter$count = 34567;
	#10 counter$count = 34568;
	#10 counter$count = 34569;
	#10 counter$count = 34570;
	#10 counter$count = 34571;
	#10 counter$count = 34572;
	#10 counter$count = 34573;
	#10 counter$count = 34574;
	#10 counter$count = 34575;
	#10 counter$count = 34576;
	#10 counter$count = 34577;
	#10 counter$count = 34578;
	#10 counter$count = 34579;
	#10 counter$count = 34580;
	#10 counter$count = 34581;
	#10 counter$count = 34582;
	#10 counter$count = 34583;
	#10 counter$count = 34584;
	#10 counter$count = 34585;
	#10 counter$count = 34586;
	#10 counter$count = 34587;
	#10 counter$count = 34588;
	#10 counter$count = 34589;
	#10 counter$count = 34590;
	#10 counter$count = 34591;
	#10 counter$count = 34592;
	#10 counter$count = 34593;
	#10 counter$count = 34594;
	#10 counter$count = 34595;
	#10 counter$count = 34596;
	#10 counter$count = 34597;
	#10 counter$count = 34598;
	#10 counter$count = 34599;
	#10 counter$count = 34600;
	#10 counter$count = 34601;
	#10 counter$count = 34602;
	#10 counter$count = 34603;
	#10 counter$count = 34604;
	#10 counter$count = 34605;
	#10 counter$count = 34606;
	#10 counter$count = 34607;
	#10 counter$count = 34608;
	#10 counter$count = 34609;
	#10 counter$count = 34610;
	#10 counter$count = 34611;
	#10 counter$count = 34612;
	#10 counter$count = 34613;
	#10 counter$count = 34614;
	#10 counter$count = 34615;
	#10 counter$count = 34616;
	#10 counter$count = 34617;
	#10 counter$count = 34618;
	#10 counter$count = 34619;
	#10 counter$count = 34620;
	#10 counter$count = 34621;
	#10 counter$count = 34622;
	#10 counter$count = 34623;
	#10 counter$count = 34624;
	#10 counter$count = 34625;
	#10 counter$count = 34626;
	#10 counter$count = 34627;
	#10 counter$count = 34628;
	#10 counter$count = 34629;
	#10 counter$count = 34630;
	#10 counter$count = 34631;
	#10 counter$count = 34632;
	#10 counter$count = 34633;
	#10 counter$count = 34634;
	#10 counter$count = 34635;
	#10 counter$count = 34636;
	#10 counter$count = 34637;
	#10 counter$count = 34638;
	#10 counter$count = 34639;
	#10 counter$count = 34640;
	#10 counter$count = 34641;
	#10 counter$count = 34642;
	#10 counter$count = 34643;
	#10 counter$count = 34644;
	#10 counter$count = 34645;
	#10 counter$count = 34646;
	#10 counter$count = 34647;
	#10 counter$count = 34648;
	#10 counter$count = 34649;
	#10 counter$count = 34650;
	#10 counter$count = 34651;
	#10 counter$count = 34652;
	#10 counter$count = 34653;
	#10 counter$count = 34654;
	#10 counter$count = 34655;
	#10 counter$count = 34656;
	#10 counter$count = 34657;
	#10 counter$count = 34658;
	#10 counter$count = 34659;
	#10 counter$count = 34660;
	#10 counter$count = 34661;
	#10 counter$count = 34662;
	#10 counter$count = 34663;
	#10 counter$count = 34664;
	#10 counter$count = 34665;
	#10 counter$count = 34666;
	#10 counter$count = 34667;
	#10 counter$count = 34668;
	#10 counter$count = 34669;
	#10 counter$count = 34670;
	#10 counter$count = 34671;
	#10 counter$count = 34672;
	#10 counter$count = 34673;
	#10 counter$count = 34674;
	#10 counter$count = 34675;
	#10 counter$count = 34676;
	#10 counter$count = 34677;
	#10 counter$count = 34678;
	#10 counter$count = 34679;
	#10 counter$count = 34680;
	#10 counter$count = 34681;
	#10 counter$count = 34682;
	#10 counter$count = 34683;
	#10 counter$count = 34684;
	#10 counter$count = 34685;
	#10 counter$count = 34686;
	#10 counter$count = 34687;
	#10 counter$count = 34688;
	#10 counter$count = 34689;
	#10 counter$count = 34690;
	#10 counter$count = 34691;
	#10 counter$count = 34692;
	#10 counter$count = 34693;
	#10 counter$count = 34694;
	#10 counter$count = 34695;
	#10 counter$count = 34696;
	#10 counter$count = 34697;
	#10 counter$count = 34698;
	#10 counter$count = 34699;
	#10 counter$count = 34700;
	#10 counter$count = 34701;
	#10 counter$count = 34702;
	#10 counter$count = 34703;
	#10 counter$count = 34704;
	#10 counter$count = 34705;
	#10 counter$count = 34706;
	#10 counter$count = 34707;
	#10 counter$count = 34708;
	#10 counter$count = 34709;
	#10 counter$count = 34710;
	#10 counter$count = 34711;
	#10 counter$count = 34712;
	#10 counter$count = 34713;
	#10 counter$count = 34714;
	#10 counter$count = 34715;
	#10 counter$count = 34716;
	#10 counter$count = 34717;
	#10 counter$count = 34718;
	#10 counter$count = 34719;
	#10 counter$count = 34720;
	#10 counter$count = 34721;
	#10 counter$count = 34722;
	#10 counter$count = 34723;
	#10 counter$count = 34724;
	#10 counter$count = 34725;
	#10 counter$count = 34726;
	#10 counter$count = 34727;
	#10 counter$count = 34728;
	#10 counter$count = 34729;
	#10 counter$count = 34730;
	#10 counter$count = 34731;
	#10 counter$count = 34732;
	#10 counter$count = 34733;
	#10 counter$count = 34734;
	#10 counter$count = 34735;
	#10 counter$count = 34736;
	#10 counter$count = 34737;
	#10 counter$count = 34738;
	#10 counter$count = 34739;
	#10 counter$count = 34740;
	#10 counter$count = 34741;
	#10 counter$count = 34742;
	#10 counter$count = 34743;
	#10 counter$count = 34744;
	#10 counter$count = 34745;
	#10 counter$count = 34746;
	#10 counter$count = 34747;
	#10 counter$count = 34748;
	#10 counter$count = 34749;
	#10 counter$count = 34750;
	#10 counter$count = 34751;
	#10 counter$count = 34752;
	#10 counter$count = 34753;
	#10 counter$count = 34754;
	#10 counter$count = 34755;
	#10 counter$count = 34756;
	#10 counter$count = 34757;
	#10 counter$count = 34758;
	#10 counter$count = 34759;
	#10 counter$count = 34760;
	#10 counter$count = 34761;
	#10 counter$count = 34762;
	#10 counter$count = 34763;
	#10 counter$count = 34764;
	#10 counter$count = 34765;
	#10 counter$count = 34766;
	#10 counter$count = 34767;
	#10 counter$count = 34768;
	#10 counter$count = 34769;
	#10 counter$count = 34770;
	#10 counter$count = 34771;
	#10 counter$count = 34772;
	#10 counter$count = 34773;
	#10 counter$count = 34774;
	#10 counter$count = 34775;
	#10 counter$count = 34776;
	#10 counter$count = 34777;
	#10 counter$count = 34778;
	#10 counter$count = 34779;
	#10 counter$count = 34780;
	#10 counter$count = 34781;
	#10 counter$count = 34782;
	#10 counter$count = 34783;
	#10 counter$count = 34784;
	#10 counter$count = 34785;
	#10 counter$count = 34786;
	#10 counter$count = 34787;
	#10 counter$count = 34788;
	#10 counter$count = 34789;
	#10 counter$count = 34790;
	#10 counter$count = 34791;
	#10 counter$count = 34792;
	#10 counter$count = 34793;
	#10 counter$count = 34794;
	#10 counter$count = 34795;
	#10 counter$count = 34796;
	#10 counter$count = 34797;
	#10 counter$count = 34798;
	#10 counter$count = 34799;
	#10 counter$count = 34800;
	#10 counter$count = 34801;
	#10 counter$count = 34802;
	#10 counter$count = 34803;
	#10 counter$count = 34804;
	#10 counter$count = 34805;
	#10 counter$count = 34806;
	#10 counter$count = 34807;
	#10 counter$count = 34808;
	#10 counter$count = 34809;
	#10 counter$count = 34810;
	#10 counter$count = 34811;
	#10 counter$count = 34812;
	#10 counter$count = 34813;
	#10 counter$count = 34814;
	#10 counter$count = 34815;
	#10 counter$count = 34816;
	#10 counter$count = 34817;
	#10 counter$count = 34818;
	#10 counter$count = 34819;
	#10 counter$count = 34820;
	#10 counter$count = 34821;
	#10 counter$count = 34822;
	#10 counter$count = 34823;
	#10 counter$count = 34824;
	#10 counter$count = 34825;
	#10 counter$count = 34826;
	#10 counter$count = 34827;
	#10 counter$count = 34828;
	#10 counter$count = 34829;
	#10 counter$count = 34830;
	#10 counter$count = 34831;
	#10 counter$count = 34832;
	#10 counter$count = 34833;
	#10 counter$count = 34834;
	#10 counter$count = 34835;
	#10 counter$count = 34836;
	#10 counter$count = 34837;
	#10 counter$count = 34838;
	#10 counter$count = 34839;
	#10 counter$count = 34840;
	#10 counter$count = 34841;
	#10 counter$count = 34842;
	#10 counter$count = 34843;
	#10 counter$count = 34844;
	#10 counter$count = 34845;
	#10 counter$count = 34846;
	#10 counter$count = 34847;
	#10 counter$count = 34848;
	#10 counter$count = 34849;
	#10 counter$count = 34850;
	#10 counter$count = 34851;
	#10 counter$count = 34852;
	#10 counter$count = 34853;
	#10 counter$count = 34854;
	#10 counter$count = 34855;
	#10 counter$count = 34856;
	#10 counter$count = 34857;
	#10 counter$count = 34858;
	#10 counter$count = 34859;
	#10 counter$count = 34860;
	#10 counter$count = 34861;
	#10 counter$count = 34862;
	#10 counter$count = 34863;
	#10 counter$count = 34864;
	#10 counter$count = 34865;
	#10 counter$count = 34866;
	#10 counter$count = 34867;
	#10 counter$count = 34868;
	#10 counter$count = 34869;
	#10 counter$count = 34870;
	#10 counter$count = 34871;
	#10 counter$count = 34872;
	#10 counter$count = 34873;
	#10 counter$count = 34874;
	#10 counter$count = 34875;
	#10 counter$count = 34876;
	#10 counter$count = 34877;
	#10 counter$count = 34878;
	#10 counter$count = 34879;
	#10 counter$count = 34880;
	#10 counter$count = 34881;
	#10 counter$count = 34882;
	#10 counter$count = 34883;
	#10 counter$count = 34884;
	#10 counter$count = 34885;
	#10 counter$count = 34886;
	#10 counter$count = 34887;
	#10 counter$count = 34888;
	#10 counter$count = 34889;
	#10 counter$count = 34890;
	#10 counter$count = 34891;
	#10 counter$count = 34892;
	#10 counter$count = 34893;
	#10 counter$count = 34894;
	#10 counter$count = 34895;
	#10 counter$count = 34896;
	#10 counter$count = 34897;
	#10 counter$count = 34898;
	#10 counter$count = 34899;
	#10 counter$count = 34900;
	#10 counter$count = 34901;
	#10 counter$count = 34902;
	#10 counter$count = 34903;
	#10 counter$count = 34904;
	#10 counter$count = 34905;
	#10 counter$count = 34906;
	#10 counter$count = 34907;
	#10 counter$count = 34908;
	#10 counter$count = 34909;
	#10 counter$count = 34910;
	#10 counter$count = 34911;
	#10 counter$count = 34912;
	#10 counter$count = 34913;
	#10 counter$count = 34914;
	#10 counter$count = 34915;
	#10 counter$count = 34916;
	#10 counter$count = 34917;
	#10 counter$count = 34918;
	#10 counter$count = 34919;
	#10 counter$count = 34920;
	#10 counter$count = 34921;
	#10 counter$count = 34922;
	#10 counter$count = 34923;
	#10 counter$count = 34924;
	#10 counter$count = 34925;
	#10 counter$count = 34926;
	#10 counter$count = 34927;
	#10 counter$count = 34928;
	#10 counter$count = 34929;
	#10 counter$count = 34930;
	#10 counter$count = 34931;
	#10 counter$count = 34932;
	#10 counter$count = 34933;
	#10 counter$count = 34934;
	#10 counter$count = 34935;
	#10 counter$count = 34936;
	#10 counter$count = 34937;
	#10 counter$count = 34938;
	#10 counter$count = 34939;
	#10 counter$count = 34940;
	#10 counter$count = 34941;
	#10 counter$count = 34942;
	#10 counter$count = 34943;
	#10 counter$count = 34944;
	#10 counter$count = 34945;
	#10 counter$count = 34946;
	#10 counter$count = 34947;
	#10 counter$count = 34948;
	#10 counter$count = 34949;
	#10 counter$count = 34950;
	#10 counter$count = 34951;
	#10 counter$count = 34952;
	#10 counter$count = 34953;
	#10 counter$count = 34954;
	#10 counter$count = 34955;
	#10 counter$count = 34956;
	#10 counter$count = 34957;
	#10 counter$count = 34958;
	#10 counter$count = 34959;
	#10 counter$count = 34960;
	#10 counter$count = 34961;
	#10 counter$count = 34962;
	#10 counter$count = 34963;
	#10 counter$count = 34964;
	#10 counter$count = 34965;
	#10 counter$count = 34966;
	#10 counter$count = 34967;
	#10 counter$count = 34968;
	#10 counter$count = 34969;
	#10 counter$count = 34970;
	#10 counter$count = 34971;
	#10 counter$count = 34972;
	#10 counter$count = 34973;
	#10 counter$count = 34974;
	#10 counter$count = 34975;
	#10 counter$count = 34976;
	#10 counter$count = 34977;
	#10 counter$count = 34978;
	#10 counter$count = 34979;
	#10 counter$count = 34980;
	#10 counter$count = 34981;
	#10 counter$count = 34982;
	#10 counter$count = 34983;
	#10 counter$count = 34984;
	#10 counter$count = 34985;
	#10 counter$count = 34986;
	#10 counter$count = 34987;
	#10 counter$count = 34988;
	#10 counter$count = 34989;
	#10 counter$count = 34990;
	#10 counter$count = 34991;
	#10 counter$count = 34992;
	#10 counter$count = 34993;
	#10 counter$count = 34994;
	#10 counter$count = 34995;
	#10 counter$count = 34996;
	#10 counter$count = 34997;
	#10 counter$count = 34998;
	#10 counter$count = 34999;
	#10 counter$count = 35000;
	#10 counter$count = 35001;
	#10 counter$count = 35002;
	#10 counter$count = 35003;
	#10 counter$count = 35004;
	#10 counter$count = 35005;
	#10 counter$count = 35006;
	#10 counter$count = 35007;
	#10 counter$count = 35008;
	#10 counter$count = 35009;
	#10 counter$count = 35010;
	#10 counter$count = 35011;
	#10 counter$count = 35012;
	#10 counter$count = 35013;
	#10 counter$count = 35014;
	#10 counter$count = 35015;
	#10 counter$count = 35016;
	#10 counter$count = 35017;
	#10 counter$count = 35018;
	#10 counter$count = 35019;
	#10 counter$count = 35020;
	#10 counter$count = 35021;
	#10 counter$count = 35022;
	#10 counter$count = 35023;
	#10 counter$count = 35024;
	#10 counter$count = 35025;
	#10 counter$count = 35026;
	#10 counter$count = 35027;
	#10 counter$count = 35028;
	#10 counter$count = 35029;
	#10 counter$count = 35030;
	#10 counter$count = 35031;
	#10 counter$count = 35032;
	#10 counter$count = 35033;
	#10 counter$count = 35034;
	#10 counter$count = 35035;
	#10 counter$count = 35036;
	#10 counter$count = 35037;
	#10 counter$count = 35038;
	#10 counter$count = 35039;
	#10 counter$count = 35040;
	#10 counter$count = 35041;
	#10 counter$count = 35042;
	#10 counter$count = 35043;
	#10 counter$count = 35044;
	#10 counter$count = 35045;
	#10 counter$count = 35046;
	#10 counter$count = 35047;
	#10 counter$count = 35048;
	#10 counter$count = 35049;
	#10 counter$count = 35050;
	#10 counter$count = 35051;
	#10 counter$count = 35052;
	#10 counter$count = 35053;
	#10 counter$count = 35054;
	#10 counter$count = 35055;
	#10 counter$count = 35056;
	#10 counter$count = 35057;
	#10 counter$count = 35058;
	#10 counter$count = 35059;
	#10 counter$count = 35060;
	#10 counter$count = 35061;
	#10 counter$count = 35062;
	#10 counter$count = 35063;
	#10 counter$count = 35064;
	#10 counter$count = 35065;
	#10 counter$count = 35066;
	#10 counter$count = 35067;
	#10 counter$count = 35068;
	#10 counter$count = 35069;
	#10 counter$count = 35070;
	#10 counter$count = 35071;
	#10 counter$count = 35072;
	#10 counter$count = 35073;
	#10 counter$count = 35074;
	#10 counter$count = 35075;
	#10 counter$count = 35076;
	#10 counter$count = 35077;
	#10 counter$count = 35078;
	#10 counter$count = 35079;
	#10 counter$count = 35080;
	#10 counter$count = 35081;
	#10 counter$count = 35082;
	#10 counter$count = 35083;
	#10 counter$count = 35084;
	#10 counter$count = 35085;
	#10 counter$count = 35086;
	#10 counter$count = 35087;
	#10 counter$count = 35088;
	#10 counter$count = 35089;
	#10 counter$count = 35090;
	#10 counter$count = 35091;
	#10 counter$count = 35092;
	#10 counter$count = 35093;
	#10 counter$count = 35094;
	#10 counter$count = 35095;
	#10 counter$count = 35096;
	#10 counter$count = 35097;
	#10 counter$count = 35098;
	#10 counter$count = 35099;
	#10 counter$count = 35100;
	#10 counter$count = 35101;
	#10 counter$count = 35102;
	#10 counter$count = 35103;
	#10 counter$count = 35104;
	#10 counter$count = 35105;
	#10 counter$count = 35106;
	#10 counter$count = 35107;
	#10 counter$count = 35108;
	#10 counter$count = 35109;
	#10 counter$count = 35110;
	#10 counter$count = 35111;
	#10 counter$count = 35112;
	#10 counter$count = 35113;
	#10 counter$count = 35114;
	#10 counter$count = 35115;
	#10 counter$count = 35116;
	#10 counter$count = 35117;
	#10 counter$count = 35118;
	#10 counter$count = 35119;
	#10 counter$count = 35120;
	#10 counter$count = 35121;
	#10 counter$count = 35122;
	#10 counter$count = 35123;
	#10 counter$count = 35124;
	#10 counter$count = 35125;
	#10 counter$count = 35126;
	#10 counter$count = 35127;
	#10 counter$count = 35128;
	#10 counter$count = 35129;
	#10 counter$count = 35130;
	#10 counter$count = 35131;
	#10 counter$count = 35132;
	#10 counter$count = 35133;
	#10 counter$count = 35134;
	#10 counter$count = 35135;
	#10 counter$count = 35136;
	#10 counter$count = 35137;
	#10 counter$count = 35138;
	#10 counter$count = 35139;
	#10 counter$count = 35140;
	#10 counter$count = 35141;
	#10 counter$count = 35142;
	#10 counter$count = 35143;
	#10 counter$count = 35144;
	#10 counter$count = 35145;
	#10 counter$count = 35146;
	#10 counter$count = 35147;
	#10 counter$count = 35148;
	#10 counter$count = 35149;
	#10 counter$count = 35150;
	#10 counter$count = 35151;
	#10 counter$count = 35152;
	#10 counter$count = 35153;
	#10 counter$count = 35154;
	#10 counter$count = 35155;
	#10 counter$count = 35156;
	#10 counter$count = 35157;
	#10 counter$count = 35158;
	#10 counter$count = 35159;
	#10 counter$count = 35160;
	#10 counter$count = 35161;
	#10 counter$count = 35162;
	#10 counter$count = 35163;
	#10 counter$count = 35164;
	#10 counter$count = 35165;
	#10 counter$count = 35166;
	#10 counter$count = 35167;
	#10 counter$count = 35168;
	#10 counter$count = 35169;
	#10 counter$count = 35170;
	#10 counter$count = 35171;
	#10 counter$count = 35172;
	#10 counter$count = 35173;
	#10 counter$count = 35174;
	#10 counter$count = 35175;
	#10 counter$count = 35176;
	#10 counter$count = 35177;
	#10 counter$count = 35178;
	#10 counter$count = 35179;
	#10 counter$count = 35180;
	#10 counter$count = 35181;
	#10 counter$count = 35182;
	#10 counter$count = 35183;
	#10 counter$count = 35184;
	#10 counter$count = 35185;
	#10 counter$count = 35186;
	#10 counter$count = 35187;
	#10 counter$count = 35188;
	#10 counter$count = 35189;
	#10 counter$count = 35190;
	#10 counter$count = 35191;
	#10 counter$count = 35192;
	#10 counter$count = 35193;
	#10 counter$count = 35194;
	#10 counter$count = 35195;
	#10 counter$count = 35196;
	#10 counter$count = 35197;
	#10 counter$count = 35198;
	#10 counter$count = 35199;
	#10 counter$count = 35200;
	#10 counter$count = 35201;
	#10 counter$count = 35202;
	#10 counter$count = 35203;
	#10 counter$count = 35204;
	#10 counter$count = 35205;
	#10 counter$count = 35206;
	#10 counter$count = 35207;
	#10 counter$count = 35208;
	#10 counter$count = 35209;
	#10 counter$count = 35210;
	#10 counter$count = 35211;
	#10 counter$count = 35212;
	#10 counter$count = 35213;
	#10 counter$count = 35214;
	#10 counter$count = 35215;
	#10 counter$count = 35216;
	#10 counter$count = 35217;
	#10 counter$count = 35218;
	#10 counter$count = 35219;
	#10 counter$count = 35220;
	#10 counter$count = 35221;
	#10 counter$count = 35222;
	#10 counter$count = 35223;
	#10 counter$count = 35224;
	#10 counter$count = 35225;
	#10 counter$count = 35226;
	#10 counter$count = 35227;
	#10 counter$count = 35228;
	#10 counter$count = 35229;
	#10 counter$count = 35230;
	#10 counter$count = 35231;
	#10 counter$count = 35232;
	#10 counter$count = 35233;
	#10 counter$count = 35234;
	#10 counter$count = 35235;
	#10 counter$count = 35236;
	#10 counter$count = 35237;
	#10 counter$count = 35238;
	#10 counter$count = 35239;
	#10 counter$count = 35240;
	#10 counter$count = 35241;
	#10 counter$count = 35242;
	#10 counter$count = 35243;
	#10 counter$count = 35244;
	#10 counter$count = 35245;
	#10 counter$count = 35246;
	#10 counter$count = 35247;
	#10 counter$count = 35248;
	#10 counter$count = 35249;
	#10 counter$count = 35250;
	#10 counter$count = 35251;
	#10 counter$count = 35252;
	#10 counter$count = 35253;
	#10 counter$count = 35254;
	#10 counter$count = 35255;
	#10 counter$count = 35256;
	#10 counter$count = 35257;
	#10 counter$count = 35258;
	#10 counter$count = 35259;
	#10 counter$count = 35260;
	#10 counter$count = 35261;
	#10 counter$count = 35262;
	#10 counter$count = 35263;
	#10 counter$count = 35264;
	#10 counter$count = 35265;
	#10 counter$count = 35266;
	#10 counter$count = 35267;
	#10 counter$count = 35268;
	#10 counter$count = 35269;
	#10 counter$count = 35270;
	#10 counter$count = 35271;
	#10 counter$count = 35272;
	#10 counter$count = 35273;
	#10 counter$count = 35274;
	#10 counter$count = 35275;
	#10 counter$count = 35276;
	#10 counter$count = 35277;
	#10 counter$count = 35278;
	#10 counter$count = 35279;
	#10 counter$count = 35280;
	#10 counter$count = 35281;
	#10 counter$count = 35282;
	#10 counter$count = 35283;
	#10 counter$count = 35284;
	#10 counter$count = 35285;
	#10 counter$count = 35286;
	#10 counter$count = 35287;
	#10 counter$count = 35288;
	#10 counter$count = 35289;
	#10 counter$count = 35290;
	#10 counter$count = 35291;
	#10 counter$count = 35292;
	#10 counter$count = 35293;
	#10 counter$count = 35294;
	#10 counter$count = 35295;
	#10 counter$count = 35296;
	#10 counter$count = 35297;
	#10 counter$count = 35298;
	#10 counter$count = 35299;
	#10 counter$count = 35300;
	#10 counter$count = 35301;
	#10 counter$count = 35302;
	#10 counter$count = 35303;
	#10 counter$count = 35304;
	#10 counter$count = 35305;
	#10 counter$count = 35306;
	#10 counter$count = 35307;
	#10 counter$count = 35308;
	#10 counter$count = 35309;
	#10 counter$count = 35310;
	#10 counter$count = 35311;
	#10 counter$count = 35312;
	#10 counter$count = 35313;
	#10 counter$count = 35314;
	#10 counter$count = 35315;
	#10 counter$count = 35316;
	#10 counter$count = 35317;
	#10 counter$count = 35318;
	#10 counter$count = 35319;
	#10 counter$count = 35320;
	#10 counter$count = 35321;
	#10 counter$count = 35322;
	#10 counter$count = 35323;
	#10 counter$count = 35324;
	#10 counter$count = 35325;
	#10 counter$count = 35326;
	#10 counter$count = 35327;
	#10 counter$count = 35328;
	#10 counter$count = 35329;
	#10 counter$count = 35330;
	#10 counter$count = 35331;
	#10 counter$count = 35332;
	#10 counter$count = 35333;
	#10 counter$count = 35334;
	#10 counter$count = 35335;
	#10 counter$count = 35336;
	#10 counter$count = 35337;
	#10 counter$count = 35338;
	#10 counter$count = 35339;
	#10 counter$count = 35340;
	#10 counter$count = 35341;
	#10 counter$count = 35342;
	#10 counter$count = 35343;
	#10 counter$count = 35344;
	#10 counter$count = 35345;
	#10 counter$count = 35346;
	#10 counter$count = 35347;
	#10 counter$count = 35348;
	#10 counter$count = 35349;
	#10 counter$count = 35350;
	#10 counter$count = 35351;
	#10 counter$count = 35352;
	#10 counter$count = 35353;
	#10 counter$count = 35354;
	#10 counter$count = 35355;
	#10 counter$count = 35356;
	#10 counter$count = 35357;
	#10 counter$count = 35358;
	#10 counter$count = 35359;
	#10 counter$count = 35360;
	#10 counter$count = 35361;
	#10 counter$count = 35362;
	#10 counter$count = 35363;
	#10 counter$count = 35364;
	#10 counter$count = 35365;
	#10 counter$count = 35366;
	#10 counter$count = 35367;
	#10 counter$count = 35368;
	#10 counter$count = 35369;
	#10 counter$count = 35370;
	#10 counter$count = 35371;
	#10 counter$count = 35372;
	#10 counter$count = 35373;
	#10 counter$count = 35374;
	#10 counter$count = 35375;
	#10 counter$count = 35376;
	#10 counter$count = 35377;
	#10 counter$count = 35378;
	#10 counter$count = 35379;
	#10 counter$count = 35380;
	#10 counter$count = 35381;
	#10 counter$count = 35382;
	#10 counter$count = 35383;
	#10 counter$count = 35384;
	#10 counter$count = 35385;
	#10 counter$count = 35386;
	#10 counter$count = 35387;
	#10 counter$count = 35388;
	#10 counter$count = 35389;
	#10 counter$count = 35390;
	#10 counter$count = 35391;
	#10 counter$count = 35392;
	#10 counter$count = 35393;
	#10 counter$count = 35394;
	#10 counter$count = 35395;
	#10 counter$count = 35396;
	#10 counter$count = 35397;
	#10 counter$count = 35398;
	#10 counter$count = 35399;
	#10 counter$count = 35400;
	#10 counter$count = 35401;
	#10 counter$count = 35402;
	#10 counter$count = 35403;
	#10 counter$count = 35404;
	#10 counter$count = 35405;
	#10 counter$count = 35406;
	#10 counter$count = 35407;
	#10 counter$count = 35408;
	#10 counter$count = 35409;
	#10 counter$count = 35410;
	#10 counter$count = 35411;
	#10 counter$count = 35412;
	#10 counter$count = 35413;
	#10 counter$count = 35414;
	#10 counter$count = 35415;
	#10 counter$count = 35416;
	#10 counter$count = 35417;
	#10 counter$count = 35418;
	#10 counter$count = 35419;
	#10 counter$count = 35420;
	#10 counter$count = 35421;
	#10 counter$count = 35422;
	#10 counter$count = 35423;
	#10 counter$count = 35424;
	#10 counter$count = 35425;
	#10 counter$count = 35426;
	#10 counter$count = 35427;
	#10 counter$count = 35428;
	#10 counter$count = 35429;
	#10 counter$count = 35430;
	#10 counter$count = 35431;
	#10 counter$count = 35432;
	#10 counter$count = 35433;
	#10 counter$count = 35434;
	#10 counter$count = 35435;
	#10 counter$count = 35436;
	#10 counter$count = 35437;
	#10 counter$count = 35438;
	#10 counter$count = 35439;
	#10 counter$count = 35440;
	#10 counter$count = 35441;
	#10 counter$count = 35442;
	#10 counter$count = 35443;
	#10 counter$count = 35444;
	#10 counter$count = 35445;
	#10 counter$count = 35446;
	#10 counter$count = 35447;
	#10 counter$count = 35448;
	#10 counter$count = 35449;
	#10 counter$count = 35450;
	#10 counter$count = 35451;
	#10 counter$count = 35452;
	#10 counter$count = 35453;
	#10 counter$count = 35454;
	#10 counter$count = 35455;
	#10 counter$count = 35456;
	#10 counter$count = 35457;
	#10 counter$count = 35458;
	#10 counter$count = 35459;
	#10 counter$count = 35460;
	#10 counter$count = 35461;
	#10 counter$count = 35462;
	#10 counter$count = 35463;
	#10 counter$count = 35464;
	#10 counter$count = 35465;
	#10 counter$count = 35466;
	#10 counter$count = 35467;
	#10 counter$count = 35468;
	#10 counter$count = 35469;
	#10 counter$count = 35470;
	#10 counter$count = 35471;
	#10 counter$count = 35472;
	#10 counter$count = 35473;
	#10 counter$count = 35474;
	#10 counter$count = 35475;
	#10 counter$count = 35476;
	#10 counter$count = 35477;
	#10 counter$count = 35478;
	#10 counter$count = 35479;
	#10 counter$count = 35480;
	#10 counter$count = 35481;
	#10 counter$count = 35482;
	#10 counter$count = 35483;
	#10 counter$count = 35484;
	#10 counter$count = 35485;
	#10 counter$count = 35486;
	#10 counter$count = 35487;
	#10 counter$count = 35488;
	#10 counter$count = 35489;
	#10 counter$count = 35490;
	#10 counter$count = 35491;
	#10 counter$count = 35492;
	#10 counter$count = 35493;
	#10 counter$count = 35494;
	#10 counter$count = 35495;
	#10 counter$count = 35496;
	#10 counter$count = 35497;
	#10 counter$count = 35498;
	#10 counter$count = 35499;
	#10 counter$count = 35500;
	#10 counter$count = 35501;
	#10 counter$count = 35502;
	#10 counter$count = 35503;
	#10 counter$count = 35504;
	#10 counter$count = 35505;
	#10 counter$count = 35506;
	#10 counter$count = 35507;
	#10 counter$count = 35508;
	#10 counter$count = 35509;
	#10 counter$count = 35510;
	#10 counter$count = 35511;
	#10 counter$count = 35512;
	#10 counter$count = 35513;
	#10 counter$count = 35514;
	#10 counter$count = 35515;
	#10 counter$count = 35516;
	#10 counter$count = 35517;
	#10 counter$count = 35518;
	#10 counter$count = 35519;
	#10 counter$count = 35520;
	#10 counter$count = 35521;
	#10 counter$count = 35522;
	#10 counter$count = 35523;
	#10 counter$count = 35524;
	#10 counter$count = 35525;
	#10 counter$count = 35526;
	#10 counter$count = 35527;
	#10 counter$count = 35528;
	#10 counter$count = 35529;
	#10 counter$count = 35530;
	#10 counter$count = 35531;
	#10 counter$count = 35532;
	#10 counter$count = 35533;
	#10 counter$count = 35534;
	#10 counter$count = 35535;
	#10 counter$count = 35536;
	#10 counter$count = 35537;
	#10 counter$count = 35538;
	#10 counter$count = 35539;
	#10 counter$count = 35540;
	#10 counter$count = 35541;
	#10 counter$count = 35542;
	#10 counter$count = 35543;
	#10 counter$count = 35544;
	#10 counter$count = 35545;
	#10 counter$count = 35546;
	#10 counter$count = 35547;
	#10 counter$count = 35548;
	#10 counter$count = 35549;
	#10 counter$count = 35550;
	#10 counter$count = 35551;
	#10 counter$count = 35552;
	#10 counter$count = 35553;
	#10 counter$count = 35554;
	#10 counter$count = 35555;
	#10 counter$count = 35556;
	#10 counter$count = 35557;
	#10 counter$count = 35558;
	#10 counter$count = 35559;
	#10 counter$count = 35560;
	#10 counter$count = 35561;
	#10 counter$count = 35562;
	#10 counter$count = 35563;
	#10 counter$count = 35564;
	#10 counter$count = 35565;
	#10 counter$count = 35566;
	#10 counter$count = 35567;
	#10 counter$count = 35568;
	#10 counter$count = 35569;
	#10 counter$count = 35570;
	#10 counter$count = 35571;
	#10 counter$count = 35572;
	#10 counter$count = 35573;
	#10 counter$count = 35574;
	#10 counter$count = 35575;
	#10 counter$count = 35576;
	#10 counter$count = 35577;
	#10 counter$count = 35578;
	#10 counter$count = 35579;
	#10 counter$count = 35580;
	#10 counter$count = 35581;
	#10 counter$count = 35582;
	#10 counter$count = 35583;
	#10 counter$count = 35584;
	#10 counter$count = 35585;
	#10 counter$count = 35586;
	#10 counter$count = 35587;
	#10 counter$count = 35588;
	#10 counter$count = 35589;
	#10 counter$count = 35590;
	#10 counter$count = 35591;
	#10 counter$count = 35592;
	#10 counter$count = 35593;
	#10 counter$count = 35594;
	#10 counter$count = 35595;
	#10 counter$count = 35596;
	#10 counter$count = 35597;
	#10 counter$count = 35598;
	#10 counter$count = 35599;
	#10 counter$count = 35600;
	#10 counter$count = 35601;
	#10 counter$count = 35602;
	#10 counter$count = 35603;
	#10 counter$count = 35604;
	#10 counter$count = 35605;
	#10 counter$count = 35606;
	#10 counter$count = 35607;
	#10 counter$count = 35608;
	#10 counter$count = 35609;
	#10 counter$count = 35610;
	#10 counter$count = 35611;
	#10 counter$count = 35612;
	#10 counter$count = 35613;
	#10 counter$count = 35614;
	#10 counter$count = 35615;
	#10 counter$count = 35616;
	#10 counter$count = 35617;
	#10 counter$count = 35618;
	#10 counter$count = 35619;
	#10 counter$count = 35620;
	#10 counter$count = 35621;
	#10 counter$count = 35622;
	#10 counter$count = 35623;
	#10 counter$count = 35624;
	#10 counter$count = 35625;
	#10 counter$count = 35626;
	#10 counter$count = 35627;
	#10 counter$count = 35628;
	#10 counter$count = 35629;
	#10 counter$count = 35630;
	#10 counter$count = 35631;
	#10 counter$count = 35632;
	#10 counter$count = 35633;
	#10 counter$count = 35634;
	#10 counter$count = 35635;
	#10 counter$count = 35636;
	#10 counter$count = 35637;
	#10 counter$count = 35638;
	#10 counter$count = 35639;
	#10 counter$count = 35640;
	#10 counter$count = 35641;
	#10 counter$count = 35642;
	#10 counter$count = 35643;
	#10 counter$count = 35644;
	#10 counter$count = 35645;
	#10 counter$count = 35646;
	#10 counter$count = 35647;
	#10 counter$count = 35648;
	#10 counter$count = 35649;
	#10 counter$count = 35650;
	#10 counter$count = 35651;
	#10 counter$count = 35652;
	#10 counter$count = 35653;
	#10 counter$count = 35654;
	#10 counter$count = 35655;
	#10 counter$count = 35656;
	#10 counter$count = 35657;
	#10 counter$count = 35658;
	#10 counter$count = 35659;
	#10 counter$count = 35660;
	#10 counter$count = 35661;
	#10 counter$count = 35662;
	#10 counter$count = 35663;
	#10 counter$count = 35664;
	#10 counter$count = 35665;
	#10 counter$count = 35666;
	#10 counter$count = 35667;
	#10 counter$count = 35668;
	#10 counter$count = 35669;
	#10 counter$count = 35670;
	#10 counter$count = 35671;
	#10 counter$count = 35672;
	#10 counter$count = 35673;
	#10 counter$count = 35674;
	#10 counter$count = 35675;
	#10 counter$count = 35676;
	#10 counter$count = 35677;
	#10 counter$count = 35678;
	#10 counter$count = 35679;
	#10 counter$count = 35680;
	#10 counter$count = 35681;
	#10 counter$count = 35682;
	#10 counter$count = 35683;
	#10 counter$count = 35684;
	#10 counter$count = 35685;
	#10 counter$count = 35686;
	#10 counter$count = 35687;
	#10 counter$count = 35688;
	#10 counter$count = 35689;
	#10 counter$count = 35690;
	#10 counter$count = 35691;
	#10 counter$count = 35692;
	#10 counter$count = 35693;
	#10 counter$count = 35694;
	#10 counter$count = 35695;
	#10 counter$count = 35696;
	#10 counter$count = 35697;
	#10 counter$count = 35698;
	#10 counter$count = 35699;
	#10 counter$count = 35700;
	#10 counter$count = 35701;
	#10 counter$count = 35702;
	#10 counter$count = 35703;
	#10 counter$count = 35704;
	#10 counter$count = 35705;
	#10 counter$count = 35706;
	#10 counter$count = 35707;
	#10 counter$count = 35708;
	#10 counter$count = 35709;
	#10 counter$count = 35710;
	#10 counter$count = 35711;
	#10 counter$count = 35712;
	#10 counter$count = 35713;
	#10 counter$count = 35714;
	#10 counter$count = 35715;
	#10 counter$count = 35716;
	#10 counter$count = 35717;
	#10 counter$count = 35718;
	#10 counter$count = 35719;
	#10 counter$count = 35720;
	#10 counter$count = 35721;
	#10 counter$count = 35722;
	#10 counter$count = 35723;
	#10 counter$count = 35724;
	#10 counter$count = 35725;
	#10 counter$count = 35726;
	#10 counter$count = 35727;
	#10 counter$count = 35728;
	#10 counter$count = 35729;
	#10 counter$count = 35730;
	#10 counter$count = 35731;
	#10 counter$count = 35732;
	#10 counter$count = 35733;
	#10 counter$count = 35734;
	#10 counter$count = 35735;
	#10 counter$count = 35736;
	#10 counter$count = 35737;
	#10 counter$count = 35738;
	#10 counter$count = 35739;
	#10 counter$count = 35740;
	#10 counter$count = 35741;
	#10 counter$count = 35742;
	#10 counter$count = 35743;
	#10 counter$count = 35744;
	#10 counter$count = 35745;
	#10 counter$count = 35746;
	#10 counter$count = 35747;
	#10 counter$count = 35748;
	#10 counter$count = 35749;
	#10 counter$count = 35750;
	#10 counter$count = 35751;
	#10 counter$count = 35752;
	#10 counter$count = 35753;
	#10 counter$count = 35754;
	#10 counter$count = 35755;
	#10 counter$count = 35756;
	#10 counter$count = 35757;
	#10 counter$count = 35758;
	#10 counter$count = 35759;
	#10 counter$count = 35760;
	#10 counter$count = 35761;
	#10 counter$count = 35762;
	#10 counter$count = 35763;
	#10 counter$count = 35764;
	#10 counter$count = 35765;
	#10 counter$count = 35766;
	#10 counter$count = 35767;
	#10 counter$count = 35768;
	#10 counter$count = 35769;
	#10 counter$count = 35770;
	#10 counter$count = 35771;
	#10 counter$count = 35772;
	#10 counter$count = 35773;
	#10 counter$count = 35774;
	#10 counter$count = 35775;
	#10 counter$count = 35776;
	#10 counter$count = 35777;
	#10 counter$count = 35778;
	#10 counter$count = 35779;
	#10 counter$count = 35780;
	#10 counter$count = 35781;
	#10 counter$count = 35782;
	#10 counter$count = 35783;
	#10 counter$count = 35784;
	#10 counter$count = 35785;
	#10 counter$count = 35786;
	#10 counter$count = 35787;
	#10 counter$count = 35788;
	#10 counter$count = 35789;
	#10 counter$count = 35790;
	#10 counter$count = 35791;
	#10 counter$count = 35792;
	#10 counter$count = 35793;
	#10 counter$count = 35794;
	#10 counter$count = 35795;
	#10 counter$count = 35796;
	#10 counter$count = 35797;
	#10 counter$count = 35798;
	#10 counter$count = 35799;
	#10 counter$count = 35800;
	#10 counter$count = 35801;
	#10 counter$count = 35802;
	#10 counter$count = 35803;
	#10 counter$count = 35804;
	#10 counter$count = 35805;
	#10 counter$count = 35806;
	#10 counter$count = 35807;
	#10 counter$count = 35808;
	#10 counter$count = 35809;
	#10 counter$count = 35810;
	#10 counter$count = 35811;
	#10 counter$count = 35812;
	#10 counter$count = 35813;
	#10 counter$count = 35814;
	#10 counter$count = 35815;
	#10 counter$count = 35816;
	#10 counter$count = 35817;
	#10 counter$count = 35818;
	#10 counter$count = 35819;
	#10 counter$count = 35820;
	#10 counter$count = 35821;
	#10 counter$count = 35822;
	#10 counter$count = 35823;
	#10 counter$count = 35824;
	#10 counter$count = 35825;
	#10 counter$count = 35826;
	#10 counter$count = 35827;
	#10 counter$count = 35828;
	#10 counter$count = 35829;
	#10 counter$count = 35830;
	#10 counter$count = 35831;
	#10 counter$count = 35832;
	#10 counter$count = 35833;
	#10 counter$count = 35834;
	#10 counter$count = 35835;
	#10 counter$count = 35836;
	#10 counter$count = 35837;
	#10 counter$count = 35838;
	#10 counter$count = 35839;
	#10 counter$count = 35840;
	#10 counter$count = 35841;
	#10 counter$count = 35842;
	#10 counter$count = 35843;
	#10 counter$count = 35844;
	#10 counter$count = 35845;
	#10 counter$count = 35846;
	#10 counter$count = 35847;
	#10 counter$count = 35848;
	#10 counter$count = 35849;
	#10 counter$count = 35850;
	#10 counter$count = 35851;
	#10 counter$count = 35852;
	#10 counter$count = 35853;
	#10 counter$count = 35854;
	#10 counter$count = 35855;
	#10 counter$count = 35856;
	#10 counter$count = 35857;
	#10 counter$count = 35858;
	#10 counter$count = 35859;
	#10 counter$count = 35860;
	#10 counter$count = 35861;
	#10 counter$count = 35862;
	#10 counter$count = 35863;
	#10 counter$count = 35864;
	#10 counter$count = 35865;
	#10 counter$count = 35866;
	#10 counter$count = 35867;
	#10 counter$count = 35868;
	#10 counter$count = 35869;
	#10 counter$count = 35870;
	#10 counter$count = 35871;
	#10 counter$count = 35872;
	#10 counter$count = 35873;
	#10 counter$count = 35874;
	#10 counter$count = 35875;
	#10 counter$count = 35876;
	#10 counter$count = 35877;
	#10 counter$count = 35878;
	#10 counter$count = 35879;
	#10 counter$count = 35880;
	#10 counter$count = 35881;
	#10 counter$count = 35882;
	#10 counter$count = 35883;
	#10 counter$count = 35884;
	#10 counter$count = 35885;
	#10 counter$count = 35886;
	#10 counter$count = 35887;
	#10 counter$count = 35888;
	#10 counter$count = 35889;
	#10 counter$count = 35890;
	#10 counter$count = 35891;
	#10 counter$count = 35892;
	#10 counter$count = 35893;
	#10 counter$count = 35894;
	#10 counter$count = 35895;
	#10 counter$count = 35896;
	#10 counter$count = 35897;
	#10 counter$count = 35898;
	#10 counter$count = 35899;
	#10 counter$count = 35900;
	#10 counter$count = 35901;
	#10 counter$count = 35902;
	#10 counter$count = 35903;
	#10 counter$count = 35904;
	#10 counter$count = 35905;
	#10 counter$count = 35906;
	#10 counter$count = 35907;
	#10 counter$count = 35908;
	#10 counter$count = 35909;
	#10 counter$count = 35910;
	#10 counter$count = 35911;
	#10 counter$count = 35912;
	#10 counter$count = 35913;
	#10 counter$count = 35914;
	#10 counter$count = 35915;
	#10 counter$count = 35916;
	#10 counter$count = 35917;
	#10 counter$count = 35918;
	#10 counter$count = 35919;
	#10 counter$count = 35920;
	#10 counter$count = 35921;
	#10 counter$count = 35922;
	#10 counter$count = 35923;
	#10 counter$count = 35924;
	#10 counter$count = 35925;
	#10 counter$count = 35926;
	#10 counter$count = 35927;
	#10 counter$count = 35928;
	#10 counter$count = 35929;
	#10 counter$count = 35930;
	#10 counter$count = 35931;
	#10 counter$count = 35932;
	#10 counter$count = 35933;
	#10 counter$count = 35934;
	#10 counter$count = 35935;
	#10 counter$count = 35936;
	#10 counter$count = 35937;
	#10 counter$count = 35938;
	#10 counter$count = 35939;
	#10 counter$count = 35940;
	#10 counter$count = 35941;
	#10 counter$count = 35942;
	#10 counter$count = 35943;
	#10 counter$count = 35944;
	#10 counter$count = 35945;
	#10 counter$count = 35946;
	#10 counter$count = 35947;
	#10 counter$count = 35948;
	#10 counter$count = 35949;
	#10 counter$count = 35950;
	#10 counter$count = 35951;
	#10 counter$count = 35952;
	#10 counter$count = 35953;
	#10 counter$count = 35954;
	#10 counter$count = 35955;
	#10 counter$count = 35956;
	#10 counter$count = 35957;
	#10 counter$count = 35958;
	#10 counter$count = 35959;
	#10 counter$count = 35960;
	#10 counter$count = 35961;
	#10 counter$count = 35962;
	#10 counter$count = 35963;
	#10 counter$count = 35964;
	#10 counter$count = 35965;
	#10 counter$count = 35966;
	#10 counter$count = 35967;
	#10 counter$count = 35968;
	#10 counter$count = 35969;
	#10 counter$count = 35970;
	#10 counter$count = 35971;
	#10 counter$count = 35972;
	#10 counter$count = 35973;
	#10 counter$count = 35974;
	#10 counter$count = 35975;
	#10 counter$count = 35976;
	#10 counter$count = 35977;
	#10 counter$count = 35978;
	#10 counter$count = 35979;
	#10 counter$count = 35980;
	#10 counter$count = 35981;
	#10 counter$count = 35982;
	#10 counter$count = 35983;
	#10 counter$count = 35984;
	#10 counter$count = 35985;
	#10 counter$count = 35986;
	#10 counter$count = 35987;
	#10 counter$count = 35988;
	#10 counter$count = 35989;
	#10 counter$count = 35990;
	#10 counter$count = 35991;
	#10 counter$count = 35992;
	#10 counter$count = 35993;
	#10 counter$count = 35994;
	#10 counter$count = 35995;
	#10 counter$count = 35996;
	#10 counter$count = 35997;
	#10 counter$count = 35998;
	#10 counter$count = 35999;
	#10 counter$count = 36000;
	#10 counter$count = 36001;
	#10 counter$count = 36002;
	#10 counter$count = 36003;
	#10 counter$count = 36004;
	#10 counter$count = 36005;
	#10 counter$count = 36006;
	#10 counter$count = 36007;
	#10 counter$count = 36008;
	#10 counter$count = 36009;
	#10 counter$count = 36010;
	#10 counter$count = 36011;
	#10 counter$count = 36012;
	#10 counter$count = 36013;
	#10 counter$count = 36014;
	#10 counter$count = 36015;
	#10 counter$count = 36016;
	#10 counter$count = 36017;
	#10 counter$count = 36018;
	#10 counter$count = 36019;
	#10 counter$count = 36020;
	#10 counter$count = 36021;
	#10 counter$count = 36022;
	#10 counter$count = 36023;
	#10 counter$count = 36024;
	#10 counter$count = 36025;
	#10 counter$count = 36026;
	#10 counter$count = 36027;
	#10 counter$count = 36028;
	#10 counter$count = 36029;
	#10 counter$count = 36030;
	#10 counter$count = 36031;
	#10 counter$count = 36032;
	#10 counter$count = 36033;
	#10 counter$count = 36034;
	#10 counter$count = 36035;
	#10 counter$count = 36036;
	#10 counter$count = 36037;
	#10 counter$count = 36038;
	#10 counter$count = 36039;
	#10 counter$count = 36040;
	#10 counter$count = 36041;
	#10 counter$count = 36042;
	#10 counter$count = 36043;
	#10 counter$count = 36044;
	#10 counter$count = 36045;
	#10 counter$count = 36046;
	#10 counter$count = 36047;
	#10 counter$count = 36048;
	#10 counter$count = 36049;
	#10 counter$count = 36050;
	#10 counter$count = 36051;
	#10 counter$count = 36052;
	#10 counter$count = 36053;
	#10 counter$count = 36054;
	#10 counter$count = 36055;
	#10 counter$count = 36056;
	#10 counter$count = 36057;
	#10 counter$count = 36058;
	#10 counter$count = 36059;
	#10 counter$count = 36060;
	#10 counter$count = 36061;
	#10 counter$count = 36062;
	#10 counter$count = 36063;
	#10 counter$count = 36064;
	#10 counter$count = 36065;
	#10 counter$count = 36066;
	#10 counter$count = 36067;
	#10 counter$count = 36068;
	#10 counter$count = 36069;
	#10 counter$count = 36070;
	#10 counter$count = 36071;
	#10 counter$count = 36072;
	#10 counter$count = 36073;
	#10 counter$count = 36074;
	#10 counter$count = 36075;
	#10 counter$count = 36076;
	#10 counter$count = 36077;
	#10 counter$count = 36078;
	#10 counter$count = 36079;
	#10 counter$count = 36080;
	#10 counter$count = 36081;
	#10 counter$count = 36082;
	#10 counter$count = 36083;
	#10 counter$count = 36084;
	#10 counter$count = 36085;
	#10 counter$count = 36086;
	#10 counter$count = 36087;
	#10 counter$count = 36088;
	#10 counter$count = 36089;
	#10 counter$count = 36090;
	#10 counter$count = 36091;
	#10 counter$count = 36092;
	#10 counter$count = 36093;
	#10 counter$count = 36094;
	#10 counter$count = 36095;
	#10 counter$count = 36096;
	#10 counter$count = 36097;
	#10 counter$count = 36098;
	#10 counter$count = 36099;
	#10 counter$count = 36100;
	#10 counter$count = 36101;
	#10 counter$count = 36102;
	#10 counter$count = 36103;
	#10 counter$count = 36104;
	#10 counter$count = 36105;
	#10 counter$count = 36106;
	#10 counter$count = 36107;
	#10 counter$count = 36108;
	#10 counter$count = 36109;
	#10 counter$count = 36110;
	#10 counter$count = 36111;
	#10 counter$count = 36112;
	#10 counter$count = 36113;
	#10 counter$count = 36114;
	#10 counter$count = 36115;
	#10 counter$count = 36116;
	#10 counter$count = 36117;
	#10 counter$count = 36118;
	#10 counter$count = 36119;
	#10 counter$count = 36120;
	#10 counter$count = 36121;
	#10 counter$count = 36122;
	#10 counter$count = 36123;
	#10 counter$count = 36124;
	#10 counter$count = 36125;
	#10 counter$count = 36126;
	#10 counter$count = 36127;
	#10 counter$count = 36128;
	#10 counter$count = 36129;
	#10 counter$count = 36130;
	#10 counter$count = 36131;
	#10 counter$count = 36132;
	#10 counter$count = 36133;
	#10 counter$count = 36134;
	#10 counter$count = 36135;
	#10 counter$count = 36136;
	#10 counter$count = 36137;
	#10 counter$count = 36138;
	#10 counter$count = 36139;
	#10 counter$count = 36140;
	#10 counter$count = 36141;
	#10 counter$count = 36142;
	#10 counter$count = 36143;
	#10 counter$count = 36144;
	#10 counter$count = 36145;
	#10 counter$count = 36146;
	#10 counter$count = 36147;
	#10 counter$count = 36148;
	#10 counter$count = 36149;
	#10 counter$count = 36150;
	#10 counter$count = 36151;
	#10 counter$count = 36152;
	#10 counter$count = 36153;
	#10 counter$count = 36154;
	#10 counter$count = 36155;
	#10 counter$count = 36156;
	#10 counter$count = 36157;
	#10 counter$count = 36158;
	#10 counter$count = 36159;
	#10 counter$count = 36160;
	#10 counter$count = 36161;
	#10 counter$count = 36162;
	#10 counter$count = 36163;
	#10 counter$count = 36164;
	#10 counter$count = 36165;
	#10 counter$count = 36166;
	#10 counter$count = 36167;
	#10 counter$count = 36168;
	#10 counter$count = 36169;
	#10 counter$count = 36170;
	#10 counter$count = 36171;
	#10 counter$count = 36172;
	#10 counter$count = 36173;
	#10 counter$count = 36174;
	#10 counter$count = 36175;
	#10 counter$count = 36176;
	#10 counter$count = 36177;
	#10 counter$count = 36178;
	#10 counter$count = 36179;
	#10 counter$count = 36180;
	#10 counter$count = 36181;
	#10 counter$count = 36182;
	#10 counter$count = 36183;
	#10 counter$count = 36184;
	#10 counter$count = 36185;
	#10 counter$count = 36186;
	#10 counter$count = 36187;
	#10 counter$count = 36188;
	#10 counter$count = 36189;
	#10 counter$count = 36190;
	#10 counter$count = 36191;
	#10 counter$count = 36192;
	#10 counter$count = 36193;
	#10 counter$count = 36194;
	#10 counter$count = 36195;
	#10 counter$count = 36196;
	#10 counter$count = 36197;
	#10 counter$count = 36198;
	#10 counter$count = 36199;
	#10 counter$count = 36200;
	#10 counter$count = 36201;
	#10 counter$count = 36202;
	#10 counter$count = 36203;
	#10 counter$count = 36204;
	#10 counter$count = 36205;
	#10 counter$count = 36206;
	#10 counter$count = 36207;
	#10 counter$count = 36208;
	#10 counter$count = 36209;
	#10 counter$count = 36210;
	#10 counter$count = 36211;
	#10 counter$count = 36212;
	#10 counter$count = 36213;
	#10 counter$count = 36214;
	#10 counter$count = 36215;
	#10 counter$count = 36216;
	#10 counter$count = 36217;
	#10 counter$count = 36218;
	#10 counter$count = 36219;
	#10 counter$count = 36220;
	#10 counter$count = 36221;
	#10 counter$count = 36222;
	#10 counter$count = 36223;
	#10 counter$count = 36224;
	#10 counter$count = 36225;
	#10 counter$count = 36226;
	#10 counter$count = 36227;
	#10 counter$count = 36228;
	#10 counter$count = 36229;
	#10 counter$count = 36230;
	#10 counter$count = 36231;
	#10 counter$count = 36232;
	#10 counter$count = 36233;
	#10 counter$count = 36234;
	#10 counter$count = 36235;
	#10 counter$count = 36236;
	#10 counter$count = 36237;
	#10 counter$count = 36238;
	#10 counter$count = 36239;
	#10 counter$count = 36240;
	#10 counter$count = 36241;
	#10 counter$count = 36242;
	#10 counter$count = 36243;
	#10 counter$count = 36244;
	#10 counter$count = 36245;
	#10 counter$count = 36246;
	#10 counter$count = 36247;
	#10 counter$count = 36248;
	#10 counter$count = 36249;
	#10 counter$count = 36250;
	#10 counter$count = 36251;
	#10 counter$count = 36252;
	#10 counter$count = 36253;
	#10 counter$count = 36254;
	#10 counter$count = 36255;
	#10 counter$count = 36256;
	#10 counter$count = 36257;
	#10 counter$count = 36258;
	#10 counter$count = 36259;
	#10 counter$count = 36260;
	#10 counter$count = 36261;
	#10 counter$count = 36262;
	#10 counter$count = 36263;
	#10 counter$count = 36264;
	#10 counter$count = 36265;
	#10 counter$count = 36266;
	#10 counter$count = 36267;
	#10 counter$count = 36268;
	#10 counter$count = 36269;
	#10 counter$count = 36270;
	#10 counter$count = 36271;
	#10 counter$count = 36272;
	#10 counter$count = 36273;
	#10 counter$count = 36274;
	#10 counter$count = 36275;
	#10 counter$count = 36276;
	#10 counter$count = 36277;
	#10 counter$count = 36278;
	#10 counter$count = 36279;
	#10 counter$count = 36280;
	#10 counter$count = 36281;
	#10 counter$count = 36282;
	#10 counter$count = 36283;
	#10 counter$count = 36284;
	#10 counter$count = 36285;
	#10 counter$count = 36286;
	#10 counter$count = 36287;
	#10 counter$count = 36288;
	#10 counter$count = 36289;
	#10 counter$count = 36290;
	#10 counter$count = 36291;
	#10 counter$count = 36292;
	#10 counter$count = 36293;
	#10 counter$count = 36294;
	#10 counter$count = 36295;
	#10 counter$count = 36296;
	#10 counter$count = 36297;
	#10 counter$count = 36298;
	#10 counter$count = 36299;
	#10 counter$count = 36300;
	#10 counter$count = 36301;
	#10 counter$count = 36302;
	#10 counter$count = 36303;
	#10 counter$count = 36304;
	#10 counter$count = 36305;
	#10 counter$count = 36306;
	#10 counter$count = 36307;
	#10 counter$count = 36308;
	#10 counter$count = 36309;
	#10 counter$count = 36310;
	#10 counter$count = 36311;
	#10 counter$count = 36312;
	#10 counter$count = 36313;
	#10 counter$count = 36314;
	#10 counter$count = 36315;
	#10 counter$count = 36316;
	#10 counter$count = 36317;
	#10 counter$count = 36318;
	#10 counter$count = 36319;
	#10 counter$count = 36320;
	#10 counter$count = 36321;
	#10 counter$count = 36322;
	#10 counter$count = 36323;
	#10 counter$count = 36324;
	#10 counter$count = 36325;
	#10 counter$count = 36326;
	#10 counter$count = 36327;
	#10 counter$count = 36328;
	#10 counter$count = 36329;
	#10 counter$count = 36330;
	#10 counter$count = 36331;
	#10 counter$count = 36332;
	#10 counter$count = 36333;
	#10 counter$count = 36334;
	#10 counter$count = 36335;
	#10 counter$count = 36336;
	#10 counter$count = 36337;
	#10 counter$count = 36338;
	#10 counter$count = 36339;
	#10 counter$count = 36340;
	#10 counter$count = 36341;
	#10 counter$count = 36342;
	#10 counter$count = 36343;
	#10 counter$count = 36344;
	#10 counter$count = 36345;
	#10 counter$count = 36346;
	#10 counter$count = 36347;
	#10 counter$count = 36348;
	#10 counter$count = 36349;
	#10 counter$count = 36350;
	#10 counter$count = 36351;
	#10 counter$count = 36352;
	#10 counter$count = 36353;
	#10 counter$count = 36354;
	#10 counter$count = 36355;
	#10 counter$count = 36356;
	#10 counter$count = 36357;
	#10 counter$count = 36358;
	#10 counter$count = 36359;
	#10 counter$count = 36360;
	#10 counter$count = 36361;
	#10 counter$count = 36362;
	#10 counter$count = 36363;
	#10 counter$count = 36364;
	#10 counter$count = 36365;
	#10 counter$count = 36366;
	#10 counter$count = 36367;
	#10 counter$count = 36368;
	#10 counter$count = 36369;
	#10 counter$count = 36370;
	#10 counter$count = 36371;
	#10 counter$count = 36372;
	#10 counter$count = 36373;
	#10 counter$count = 36374;
	#10 counter$count = 36375;
	#10 counter$count = 36376;
	#10 counter$count = 36377;
	#10 counter$count = 36378;
	#10 counter$count = 36379;
	#10 counter$count = 36380;
	#10 counter$count = 36381;
	#10 counter$count = 36382;
	#10 counter$count = 36383;
	#10 counter$count = 36384;
	#10 counter$count = 36385;
	#10 counter$count = 36386;
	#10 counter$count = 36387;
	#10 counter$count = 36388;
	#10 counter$count = 36389;
	#10 counter$count = 36390;
	#10 counter$count = 36391;
	#10 counter$count = 36392;
	#10 counter$count = 36393;
	#10 counter$count = 36394;
	#10 counter$count = 36395;
	#10 counter$count = 36396;
	#10 counter$count = 36397;
	#10 counter$count = 36398;
	#10 counter$count = 36399;
	#10 counter$count = 36400;
	#10 counter$count = 36401;
	#10 counter$count = 36402;
	#10 counter$count = 36403;
	#10 counter$count = 36404;
	#10 counter$count = 36405;
	#10 counter$count = 36406;
	#10 counter$count = 36407;
	#10 counter$count = 36408;
	#10 counter$count = 36409;
	#10 counter$count = 36410;
	#10 counter$count = 36411;
	#10 counter$count = 36412;
	#10 counter$count = 36413;
	#10 counter$count = 36414;
	#10 counter$count = 36415;
	#10 counter$count = 36416;
	#10 counter$count = 36417;
	#10 counter$count = 36418;
	#10 counter$count = 36419;
	#10 counter$count = 36420;
	#10 counter$count = 36421;
	#10 counter$count = 36422;
	#10 counter$count = 36423;
	#10 counter$count = 36424;
	#10 counter$count = 36425;
	#10 counter$count = 36426;
	#10 counter$count = 36427;
	#10 counter$count = 36428;
	#10 counter$count = 36429;
	#10 counter$count = 36430;
	#10 counter$count = 36431;
	#10 counter$count = 36432;
	#10 counter$count = 36433;
	#10 counter$count = 36434;
	#10 counter$count = 36435;
	#10 counter$count = 36436;
	#10 counter$count = 36437;
	#10 counter$count = 36438;
	#10 counter$count = 36439;
	#10 counter$count = 36440;
	#10 counter$count = 36441;
	#10 counter$count = 36442;
	#10 counter$count = 36443;
	#10 counter$count = 36444;
	#10 counter$count = 36445;
	#10 counter$count = 36446;
	#10 counter$count = 36447;
	#10 counter$count = 36448;
	#10 counter$count = 36449;
	#10 counter$count = 36450;
	#10 counter$count = 36451;
	#10 counter$count = 36452;
	#10 counter$count = 36453;
	#10 counter$count = 36454;
	#10 counter$count = 36455;
	#10 counter$count = 36456;
	#10 counter$count = 36457;
	#10 counter$count = 36458;
	#10 counter$count = 36459;
	#10 counter$count = 36460;
	#10 counter$count = 36461;
	#10 counter$count = 36462;
	#10 counter$count = 36463;
	#10 counter$count = 36464;
	#10 counter$count = 36465;
	#10 counter$count = 36466;
	#10 counter$count = 36467;
	#10 counter$count = 36468;
	#10 counter$count = 36469;
	#10 counter$count = 36470;
	#10 counter$count = 36471;
	#10 counter$count = 36472;
	#10 counter$count = 36473;
	#10 counter$count = 36474;
	#10 counter$count = 36475;
	#10 counter$count = 36476;
	#10 counter$count = 36477;
	#10 counter$count = 36478;
	#10 counter$count = 36479;
	#10 counter$count = 36480;
	#10 counter$count = 36481;
	#10 counter$count = 36482;
	#10 counter$count = 36483;
	#10 counter$count = 36484;
	#10 counter$count = 36485;
	#10 counter$count = 36486;
	#10 counter$count = 36487;
	#10 counter$count = 36488;
	#10 counter$count = 36489;
	#10 counter$count = 36490;
	#10 counter$count = 36491;
	#10 counter$count = 36492;
	#10 counter$count = 36493;
	#10 counter$count = 36494;
	#10 counter$count = 36495;
	#10 counter$count = 36496;
	#10 counter$count = 36497;
	#10 counter$count = 36498;
	#10 counter$count = 36499;
	#10 counter$count = 36500;
	#10 counter$count = 36501;
	#10 counter$count = 36502;
	#10 counter$count = 36503;
	#10 counter$count = 36504;
	#10 counter$count = 36505;
	#10 counter$count = 36506;
	#10 counter$count = 36507;
	#10 counter$count = 36508;
	#10 counter$count = 36509;
	#10 counter$count = 36510;
	#10 counter$count = 36511;
	#10 counter$count = 36512;
	#10 counter$count = 36513;
	#10 counter$count = 36514;
	#10 counter$count = 36515;
	#10 counter$count = 36516;
	#10 counter$count = 36517;
	#10 counter$count = 36518;
	#10 counter$count = 36519;
	#10 counter$count = 36520;
	#10 counter$count = 36521;
	#10 counter$count = 36522;
	#10 counter$count = 36523;
	#10 counter$count = 36524;
	#10 counter$count = 36525;
	#10 counter$count = 36526;
	#10 counter$count = 36527;
	#10 counter$count = 36528;
	#10 counter$count = 36529;
	#10 counter$count = 36530;
	#10 counter$count = 36531;
	#10 counter$count = 36532;
	#10 counter$count = 36533;
	#10 counter$count = 36534;
	#10 counter$count = 36535;
	#10 counter$count = 36536;
	#10 counter$count = 36537;
	#10 counter$count = 36538;
	#10 counter$count = 36539;
	#10 counter$count = 36540;
	#10 counter$count = 36541;
	#10 counter$count = 36542;
	#10 counter$count = 36543;
	#10 counter$count = 36544;
	#10 counter$count = 36545;
	#10 counter$count = 36546;
	#10 counter$count = 36547;
	#10 counter$count = 36548;
	#10 counter$count = 36549;
	#10 counter$count = 36550;
	#10 counter$count = 36551;
	#10 counter$count = 36552;
	#10 counter$count = 36553;
	#10 counter$count = 36554;
	#10 counter$count = 36555;
	#10 counter$count = 36556;
	#10 counter$count = 36557;
	#10 counter$count = 36558;
	#10 counter$count = 36559;
	#10 counter$count = 36560;
	#10 counter$count = 36561;
	#10 counter$count = 36562;
	#10 counter$count = 36563;
	#10 counter$count = 36564;
	#10 counter$count = 36565;
	#10 counter$count = 36566;
	#10 counter$count = 36567;
	#10 counter$count = 36568;
	#10 counter$count = 36569;
	#10 counter$count = 36570;
	#10 counter$count = 36571;
	#10 counter$count = 36572;
	#10 counter$count = 36573;
	#10 counter$count = 36574;
	#10 counter$count = 36575;
	#10 counter$count = 36576;
	#10 counter$count = 36577;
	#10 counter$count = 36578;
	#10 counter$count = 36579;
	#10 counter$count = 36580;
	#10 counter$count = 36581;
	#10 counter$count = 36582;
	#10 counter$count = 36583;
	#10 counter$count = 36584;
	#10 counter$count = 36585;
	#10 counter$count = 36586;
	#10 counter$count = 36587;
	#10 counter$count = 36588;
	#10 counter$count = 36589;
	#10 counter$count = 36590;
	#10 counter$count = 36591;
	#10 counter$count = 36592;
	#10 counter$count = 36593;
	#10 counter$count = 36594;
	#10 counter$count = 36595;
	#10 counter$count = 36596;
	#10 counter$count = 36597;
	#10 counter$count = 36598;
	#10 counter$count = 36599;
	#10 counter$count = 36600;
	#10 counter$count = 36601;
	#10 counter$count = 36602;
	#10 counter$count = 36603;
	#10 counter$count = 36604;
	#10 counter$count = 36605;
	#10 counter$count = 36606;
	#10 counter$count = 36607;
	#10 counter$count = 36608;
	#10 counter$count = 36609;
	#10 counter$count = 36610;
	#10 counter$count = 36611;
	#10 counter$count = 36612;
	#10 counter$count = 36613;
	#10 counter$count = 36614;
	#10 counter$count = 36615;
	#10 counter$count = 36616;
	#10 counter$count = 36617;
	#10 counter$count = 36618;
	#10 counter$count = 36619;
	#10 counter$count = 36620;
	#10 counter$count = 36621;
	#10 counter$count = 36622;
	#10 counter$count = 36623;
	#10 counter$count = 36624;
	#10 counter$count = 36625;
	#10 counter$count = 36626;
	#10 counter$count = 36627;
	#10 counter$count = 36628;
	#10 counter$count = 36629;
	#10 counter$count = 36630;
	#10 counter$count = 36631;
	#10 counter$count = 36632;
	#10 counter$count = 36633;
	#10 counter$count = 36634;
	#10 counter$count = 36635;
	#10 counter$count = 36636;
	#10 counter$count = 36637;
	#10 counter$count = 36638;
	#10 counter$count = 36639;
	#10 counter$count = 36640;
	#10 counter$count = 36641;
	#10 counter$count = 36642;
	#10 counter$count = 36643;
	#10 counter$count = 36644;
	#10 counter$count = 36645;
	#10 counter$count = 36646;
	#10 counter$count = 36647;
	#10 counter$count = 36648;
	#10 counter$count = 36649;
	#10 counter$count = 36650;
	#10 counter$count = 36651;
	#10 counter$count = 36652;
	#10 counter$count = 36653;
	#10 counter$count = 36654;
	#10 counter$count = 36655;
	#10 counter$count = 36656;
	#10 counter$count = 36657;
	#10 counter$count = 36658;
	#10 counter$count = 36659;
	#10 counter$count = 36660;
	#10 counter$count = 36661;
	#10 counter$count = 36662;
	#10 counter$count = 36663;
	#10 counter$count = 36664;
	#10 counter$count = 36665;
	#10 counter$count = 36666;
	#10 counter$count = 36667;
	#10 counter$count = 36668;
	#10 counter$count = 36669;
	#10 counter$count = 36670;
	#10 counter$count = 36671;
	#10 counter$count = 36672;
	#10 counter$count = 36673;
	#10 counter$count = 36674;
	#10 counter$count = 36675;
	#10 counter$count = 36676;
	#10 counter$count = 36677;
	#10 counter$count = 36678;
	#10 counter$count = 36679;
	#10 counter$count = 36680;
	#10 counter$count = 36681;
	#10 counter$count = 36682;
	#10 counter$count = 36683;
	#10 counter$count = 36684;
	#10 counter$count = 36685;
	#10 counter$count = 36686;
	#10 counter$count = 36687;
	#10 counter$count = 36688;
	#10 counter$count = 36689;
	#10 counter$count = 36690;
	#10 counter$count = 36691;
	#10 counter$count = 36692;
	#10 counter$count = 36693;
	#10 counter$count = 36694;
	#10 counter$count = 36695;
	#10 counter$count = 36696;
	#10 counter$count = 36697;
	#10 counter$count = 36698;
	#10 counter$count = 36699;
	#10 counter$count = 36700;
	#10 counter$count = 36701;
	#10 counter$count = 36702;
	#10 counter$count = 36703;
	#10 counter$count = 36704;
	#10 counter$count = 36705;
	#10 counter$count = 36706;
	#10 counter$count = 36707;
	#10 counter$count = 36708;
	#10 counter$count = 36709;
	#10 counter$count = 36710;
	#10 counter$count = 36711;
	#10 counter$count = 36712;
	#10 counter$count = 36713;
	#10 counter$count = 36714;
	#10 counter$count = 36715;
	#10 counter$count = 36716;
	#10 counter$count = 36717;
	#10 counter$count = 36718;
	#10 counter$count = 36719;
	#10 counter$count = 36720;
	#10 counter$count = 36721;
	#10 counter$count = 36722;
	#10 counter$count = 36723;
	#10 counter$count = 36724;
	#10 counter$count = 36725;
	#10 counter$count = 36726;
	#10 counter$count = 36727;
	#10 counter$count = 36728;
	#10 counter$count = 36729;
	#10 counter$count = 36730;
	#10 counter$count = 36731;
	#10 counter$count = 36732;
	#10 counter$count = 36733;
	#10 counter$count = 36734;
	#10 counter$count = 36735;
	#10 counter$count = 36736;
	#10 counter$count = 36737;
	#10 counter$count = 36738;
	#10 counter$count = 36739;
	#10 counter$count = 36740;
	#10 counter$count = 36741;
	#10 counter$count = 36742;
	#10 counter$count = 36743;
	#10 counter$count = 36744;
	#10 counter$count = 36745;
	#10 counter$count = 36746;
	#10 counter$count = 36747;
	#10 counter$count = 36748;
	#10 counter$count = 36749;
	#10 counter$count = 36750;
	#10 counter$count = 36751;
	#10 counter$count = 36752;
	#10 counter$count = 36753;
	#10 counter$count = 36754;
	#10 counter$count = 36755;
	#10 counter$count = 36756;
	#10 counter$count = 36757;
	#10 counter$count = 36758;
	#10 counter$count = 36759;
	#10 counter$count = 36760;
	#10 counter$count = 36761;
	#10 counter$count = 36762;
	#10 counter$count = 36763;
	#10 counter$count = 36764;
	#10 counter$count = 36765;
	#10 counter$count = 36766;
	#10 counter$count = 36767;
	#10 counter$count = 36768;
	#10 counter$count = 36769;
	#10 counter$count = 36770;
	#10 counter$count = 36771;
	#10 counter$count = 36772;
	#10 counter$count = 36773;
	#10 counter$count = 36774;
	#10 counter$count = 36775;
	#10 counter$count = 36776;
	#10 counter$count = 36777;
	#10 counter$count = 36778;
	#10 counter$count = 36779;
	#10 counter$count = 36780;
	#10 counter$count = 36781;
	#10 counter$count = 36782;
	#10 counter$count = 36783;
	#10 counter$count = 36784;
	#10 counter$count = 36785;
	#10 counter$count = 36786;
	#10 counter$count = 36787;
	#10 counter$count = 36788;
	#10 counter$count = 36789;
	#10 counter$count = 36790;
	#10 counter$count = 36791;
	#10 counter$count = 36792;
	#10 counter$count = 36793;
	#10 counter$count = 36794;
	#10 counter$count = 36795;
	#10 counter$count = 36796;
	#10 counter$count = 36797;
	#10 counter$count = 36798;
	#10 counter$count = 36799;
	#10 counter$count = 36800;
	#10 counter$count = 36801;
	#10 counter$count = 36802;
	#10 counter$count = 36803;
	#10 counter$count = 36804;
	#10 counter$count = 36805;
	#10 counter$count = 36806;
	#10 counter$count = 36807;
	#10 counter$count = 36808;
	#10 counter$count = 36809;
	#10 counter$count = 36810;
	#10 counter$count = 36811;
	#10 counter$count = 36812;
	#10 counter$count = 36813;
	#10 counter$count = 36814;
	#10 counter$count = 36815;
	#10 counter$count = 36816;
	#10 counter$count = 36817;
	#10 counter$count = 36818;
	#10 counter$count = 36819;
	#10 counter$count = 36820;
	#10 counter$count = 36821;
	#10 counter$count = 36822;
	#10 counter$count = 36823;
	#10 counter$count = 36824;
	#10 counter$count = 36825;
	#10 counter$count = 36826;
	#10 counter$count = 36827;
	#10 counter$count = 36828;
	#10 counter$count = 36829;
	#10 counter$count = 36830;
	#10 counter$count = 36831;
	#10 counter$count = 36832;
	#10 counter$count = 36833;
	#10 counter$count = 36834;
	#10 counter$count = 36835;
	#10 counter$count = 36836;
	#10 counter$count = 36837;
	#10 counter$count = 36838;
	#10 counter$count = 36839;
	#10 counter$count = 36840;
	#10 counter$count = 36841;
	#10 counter$count = 36842;
	#10 counter$count = 36843;
	#10 counter$count = 36844;
	#10 counter$count = 36845;
	#10 counter$count = 36846;
	#10 counter$count = 36847;
	#10 counter$count = 36848;
	#10 counter$count = 36849;
	#10 counter$count = 36850;
	#10 counter$count = 36851;
	#10 counter$count = 36852;
	#10 counter$count = 36853;
	#10 counter$count = 36854;
	#10 counter$count = 36855;
	#10 counter$count = 36856;
	#10 counter$count = 36857;
	#10 counter$count = 36858;
	#10 counter$count = 36859;
	#10 counter$count = 36860;
	#10 counter$count = 36861;
	#10 counter$count = 36862;
	#10 counter$count = 36863;
	#10 counter$count = 36864;
	#10 counter$count = 36865;
	#10 counter$count = 36866;
	#10 counter$count = 36867;
	#10 counter$count = 36868;
	#10 counter$count = 36869;
	#10 counter$count = 36870;
	#10 counter$count = 36871;
	#10 counter$count = 36872;
	#10 counter$count = 36873;
	#10 counter$count = 36874;
	#10 counter$count = 36875;
	#10 counter$count = 36876;
	#10 counter$count = 36877;
	#10 counter$count = 36878;
	#10 counter$count = 36879;
	#10 counter$count = 36880;
	#10 counter$count = 36881;
	#10 counter$count = 36882;
	#10 counter$count = 36883;
	#10 counter$count = 36884;
	#10 counter$count = 36885;
	#10 counter$count = 36886;
	#10 counter$count = 36887;
	#10 counter$count = 36888;
	#10 counter$count = 36889;
	#10 counter$count = 36890;
	#10 counter$count = 36891;
	#10 counter$count = 36892;
	#10 counter$count = 36893;
	#10 counter$count = 36894;
	#10 counter$count = 36895;
	#10 counter$count = 36896;
	#10 counter$count = 36897;
	#10 counter$count = 36898;
	#10 counter$count = 36899;
	#10 counter$count = 36900;
	#10 counter$count = 36901;
	#10 counter$count = 36902;
	#10 counter$count = 36903;
	#10 counter$count = 36904;
	#10 counter$count = 36905;
	#10 counter$count = 36906;
	#10 counter$count = 36907;
	#10 counter$count = 36908;
	#10 counter$count = 36909;
	#10 counter$count = 36910;
	#10 counter$count = 36911;
	#10 counter$count = 36912;
	#10 counter$count = 36913;
	#10 counter$count = 36914;
	#10 counter$count = 36915;
	#10 counter$count = 36916;
	#10 counter$count = 36917;
	#10 counter$count = 36918;
	#10 counter$count = 36919;
	#10 counter$count = 36920;
	#10 counter$count = 36921;
	#10 counter$count = 36922;
	#10 counter$count = 36923;
	#10 counter$count = 36924;
	#10 counter$count = 36925;
	#10 counter$count = 36926;
	#10 counter$count = 36927;
	#10 counter$count = 36928;
	#10 counter$count = 36929;
	#10 counter$count = 36930;
	#10 counter$count = 36931;
	#10 counter$count = 36932;
	#10 counter$count = 36933;
	#10 counter$count = 36934;
	#10 counter$count = 36935;
	#10 counter$count = 36936;
	#10 counter$count = 36937;
	#10 counter$count = 36938;
	#10 counter$count = 36939;
	#10 counter$count = 36940;
	#10 counter$count = 36941;
	#10 counter$count = 36942;
	#10 counter$count = 36943;
	#10 counter$count = 36944;
	#10 counter$count = 36945;
	#10 counter$count = 36946;
	#10 counter$count = 36947;
	#10 counter$count = 36948;
	#10 counter$count = 36949;
	#10 counter$count = 36950;
	#10 counter$count = 36951;
	#10 counter$count = 36952;
	#10 counter$count = 36953;
	#10 counter$count = 36954;
	#10 counter$count = 36955;
	#10 counter$count = 36956;
	#10 counter$count = 36957;
	#10 counter$count = 36958;
	#10 counter$count = 36959;
	#10 counter$count = 36960;
	#10 counter$count = 36961;
	#10 counter$count = 36962;
	#10 counter$count = 36963;
	#10 counter$count = 36964;
	#10 counter$count = 36965;
	#10 counter$count = 36966;
	#10 counter$count = 36967;
	#10 counter$count = 36968;
	#10 counter$count = 36969;
	#10 counter$count = 36970;
	#10 counter$count = 36971;
	#10 counter$count = 36972;
	#10 counter$count = 36973;
	#10 counter$count = 36974;
	#10 counter$count = 36975;
	#10 counter$count = 36976;
	#10 counter$count = 36977;
	#10 counter$count = 36978;
	#10 counter$count = 36979;
	#10 counter$count = 36980;
	#10 counter$count = 36981;
	#10 counter$count = 36982;
	#10 counter$count = 36983;
	#10 counter$count = 36984;
	#10 counter$count = 36985;
	#10 counter$count = 36986;
	#10 counter$count = 36987;
	#10 counter$count = 36988;
	#10 counter$count = 36989;
	#10 counter$count = 36990;
	#10 counter$count = 36991;
	#10 counter$count = 36992;
	#10 counter$count = 36993;
	#10 counter$count = 36994;
	#10 counter$count = 36995;
	#10 counter$count = 36996;
	#10 counter$count = 36997;
	#10 counter$count = 36998;
	#10 counter$count = 36999;
	#10 counter$count = 37000;
	#10 counter$count = 37001;
	#10 counter$count = 37002;
	#10 counter$count = 37003;
	#10 counter$count = 37004;
	#10 counter$count = 37005;
	#10 counter$count = 37006;
	#10 counter$count = 37007;
	#10 counter$count = 37008;
	#10 counter$count = 37009;
	#10 counter$count = 37010;
	#10 counter$count = 37011;
	#10 counter$count = 37012;
	#10 counter$count = 37013;
	#10 counter$count = 37014;
	#10 counter$count = 37015;
	#10 counter$count = 37016;
	#10 counter$count = 37017;
	#10 counter$count = 37018;
	#10 counter$count = 37019;
	#10 counter$count = 37020;
	#10 counter$count = 37021;
	#10 counter$count = 37022;
	#10 counter$count = 37023;
	#10 counter$count = 37024;
	#10 counter$count = 37025;
	#10 counter$count = 37026;
	#10 counter$count = 37027;
	#10 counter$count = 37028;
	#10 counter$count = 37029;
	#10 counter$count = 37030;
	#10 counter$count = 37031;
	#10 counter$count = 37032;
	#10 counter$count = 37033;
	#10 counter$count = 37034;
	#10 counter$count = 37035;
	#10 counter$count = 37036;
	#10 counter$count = 37037;
	#10 counter$count = 37038;
	#10 counter$count = 37039;
	#10 counter$count = 37040;
	#10 counter$count = 37041;
	#10 counter$count = 37042;
	#10 counter$count = 37043;
	#10 counter$count = 37044;
	#10 counter$count = 37045;
	#10 counter$count = 37046;
	#10 counter$count = 37047;
	#10 counter$count = 37048;
	#10 counter$count = 37049;
	#10 counter$count = 37050;
	#10 counter$count = 37051;
	#10 counter$count = 37052;
	#10 counter$count = 37053;
	#10 counter$count = 37054;
	#10 counter$count = 37055;
	#10 counter$count = 37056;
	#10 counter$count = 37057;
	#10 counter$count = 37058;
	#10 counter$count = 37059;
	#10 counter$count = 37060;
	#10 counter$count = 37061;
	#10 counter$count = 37062;
	#10 counter$count = 37063;
	#10 counter$count = 37064;
	#10 counter$count = 37065;
	#10 counter$count = 37066;
	#10 counter$count = 37067;
	#10 counter$count = 37068;
	#10 counter$count = 37069;
	#10 counter$count = 37070;
	#10 counter$count = 37071;
	#10 counter$count = 37072;
	#10 counter$count = 37073;
	#10 counter$count = 37074;
	#10 counter$count = 37075;
	#10 counter$count = 37076;
	#10 counter$count = 37077;
	#10 counter$count = 37078;
	#10 counter$count = 37079;
	#10 counter$count = 37080;
	#10 counter$count = 37081;
	#10 counter$count = 37082;
	#10 counter$count = 37083;
	#10 counter$count = 37084;
	#10 counter$count = 37085;
	#10 counter$count = 37086;
	#10 counter$count = 37087;
	#10 counter$count = 37088;
	#10 counter$count = 37089;
	#10 counter$count = 37090;
	#10 counter$count = 37091;
	#10 counter$count = 37092;
	#10 counter$count = 37093;
	#10 counter$count = 37094;
	#10 counter$count = 37095;
	#10 counter$count = 37096;
	#10 counter$count = 37097;
	#10 counter$count = 37098;
	#10 counter$count = 37099;
	#10 counter$count = 37100;
	#10 counter$count = 37101;
	#10 counter$count = 37102;
	#10 counter$count = 37103;
	#10 counter$count = 37104;
	#10 counter$count = 37105;
	#10 counter$count = 37106;
	#10 counter$count = 37107;
	#10 counter$count = 37108;
	#10 counter$count = 37109;
	#10 counter$count = 37110;
	#10 counter$count = 37111;
	#10 counter$count = 37112;
	#10 counter$count = 37113;
	#10 counter$count = 37114;
	#10 counter$count = 37115;
	#10 counter$count = 37116;
	#10 counter$count = 37117;
	#10 counter$count = 37118;
	#10 counter$count = 37119;
	#10 counter$count = 37120;
	#10 counter$count = 37121;
	#10 counter$count = 37122;
	#10 counter$count = 37123;
	#10 counter$count = 37124;
	#10 counter$count = 37125;
	#10 counter$count = 37126;
	#10 counter$count = 37127;
	#10 counter$count = 37128;
	#10 counter$count = 37129;
	#10 counter$count = 37130;
	#10 counter$count = 37131;
	#10 counter$count = 37132;
	#10 counter$count = 37133;
	#10 counter$count = 37134;
	#10 counter$count = 37135;
	#10 counter$count = 37136;
	#10 counter$count = 37137;
	#10 counter$count = 37138;
	#10 counter$count = 37139;
	#10 counter$count = 37140;
	#10 counter$count = 37141;
	#10 counter$count = 37142;
	#10 counter$count = 37143;
	#10 counter$count = 37144;
	#10 counter$count = 37145;
	#10 counter$count = 37146;
	#10 counter$count = 37147;
	#10 counter$count = 37148;
	#10 counter$count = 37149;
	#10 counter$count = 37150;
	#10 counter$count = 37151;
	#10 counter$count = 37152;
	#10 counter$count = 37153;
	#10 counter$count = 37154;
	#10 counter$count = 37155;
	#10 counter$count = 37156;
	#10 counter$count = 37157;
	#10 counter$count = 37158;
	#10 counter$count = 37159;
	#10 counter$count = 37160;
	#10 counter$count = 37161;
	#10 counter$count = 37162;
	#10 counter$count = 37163;
	#10 counter$count = 37164;
	#10 counter$count = 37165;
	#10 counter$count = 37166;
	#10 counter$count = 37167;
	#10 counter$count = 37168;
	#10 counter$count = 37169;
	#10 counter$count = 37170;
	#10 counter$count = 37171;
	#10 counter$count = 37172;
	#10 counter$count = 37173;
	#10 counter$count = 37174;
	#10 counter$count = 37175;
	#10 counter$count = 37176;
	#10 counter$count = 37177;
	#10 counter$count = 37178;
	#10 counter$count = 37179;
	#10 counter$count = 37180;
	#10 counter$count = 37181;
	#10 counter$count = 37182;
	#10 counter$count = 37183;
	#10 counter$count = 37184;
	#10 counter$count = 37185;
	#10 counter$count = 37186;
	#10 counter$count = 37187;
	#10 counter$count = 37188;
	#10 counter$count = 37189;
	#10 counter$count = 37190;
	#10 counter$count = 37191;
	#10 counter$count = 37192;
	#10 counter$count = 37193;
	#10 counter$count = 37194;
	#10 counter$count = 37195;
	#10 counter$count = 37196;
	#10 counter$count = 37197;
	#10 counter$count = 37198;
	#10 counter$count = 37199;
	#10 counter$count = 37200;
	#10 counter$count = 37201;
	#10 counter$count = 37202;
	#10 counter$count = 37203;
	#10 counter$count = 37204;
	#10 counter$count = 37205;
	#10 counter$count = 37206;
	#10 counter$count = 37207;
	#10 counter$count = 37208;
	#10 counter$count = 37209;
	#10 counter$count = 37210;
	#10 counter$count = 37211;
	#10 counter$count = 37212;
	#10 counter$count = 37213;
	#10 counter$count = 37214;
	#10 counter$count = 37215;
	#10 counter$count = 37216;
	#10 counter$count = 37217;
	#10 counter$count = 37218;
	#10 counter$count = 37219;
	#10 counter$count = 37220;
	#10 counter$count = 37221;
	#10 counter$count = 37222;
	#10 counter$count = 37223;
	#10 counter$count = 37224;
	#10 counter$count = 37225;
	#10 counter$count = 37226;
	#10 counter$count = 37227;
	#10 counter$count = 37228;
	#10 counter$count = 37229;
	#10 counter$count = 37230;
	#10 counter$count = 37231;
	#10 counter$count = 37232;
	#10 counter$count = 37233;
	#10 counter$count = 37234;
	#10 counter$count = 37235;
	#10 counter$count = 37236;
	#10 counter$count = 37237;
	#10 counter$count = 37238;
	#10 counter$count = 37239;
	#10 counter$count = 37240;
	#10 counter$count = 37241;
	#10 counter$count = 37242;
	#10 counter$count = 37243;
	#10 counter$count = 37244;
	#10 counter$count = 37245;
	#10 counter$count = 37246;
	#10 counter$count = 37247;
	#10 counter$count = 37248;
	#10 counter$count = 37249;
	#10 counter$count = 37250;
	#10 counter$count = 37251;
	#10 counter$count = 37252;
	#10 counter$count = 37253;
	#10 counter$count = 37254;
	#10 counter$count = 37255;
	#10 counter$count = 37256;
	#10 counter$count = 37257;
	#10 counter$count = 37258;
	#10 counter$count = 37259;
	#10 counter$count = 37260;
	#10 counter$count = 37261;
	#10 counter$count = 37262;
	#10 counter$count = 37263;
	#10 counter$count = 37264;
	#10 counter$count = 37265;
	#10 counter$count = 37266;
	#10 counter$count = 37267;
	#10 counter$count = 37268;
	#10 counter$count = 37269;
	#10 counter$count = 37270;
	#10 counter$count = 37271;
	#10 counter$count = 37272;
	#10 counter$count = 37273;
	#10 counter$count = 37274;
	#10 counter$count = 37275;
	#10 counter$count = 37276;
	#10 counter$count = 37277;
	#10 counter$count = 37278;
	#10 counter$count = 37279;
	#10 counter$count = 37280;
	#10 counter$count = 37281;
	#10 counter$count = 37282;
	#10 counter$count = 37283;
	#10 counter$count = 37284;
	#10 counter$count = 37285;
	#10 counter$count = 37286;
	#10 counter$count = 37287;
	#10 counter$count = 37288;
	#10 counter$count = 37289;
	#10 counter$count = 37290;
	#10 counter$count = 37291;
	#10 counter$count = 37292;
	#10 counter$count = 37293;
	#10 counter$count = 37294;
	#10 counter$count = 37295;
	#10 counter$count = 37296;
	#10 counter$count = 37297;
	#10 counter$count = 37298;
	#10 counter$count = 37299;
	#10 counter$count = 37300;
	#10 counter$count = 37301;
	#10 counter$count = 37302;
	#10 counter$count = 37303;
	#10 counter$count = 37304;
	#10 counter$count = 37305;
	#10 counter$count = 37306;
	#10 counter$count = 37307;
	#10 counter$count = 37308;
	#10 counter$count = 37309;
	#10 counter$count = 37310;
	#10 counter$count = 37311;
	#10 counter$count = 37312;
	#10 counter$count = 37313;
	#10 counter$count = 37314;
	#10 counter$count = 37315;
	#10 counter$count = 37316;
	#10 counter$count = 37317;
	#10 counter$count = 37318;
	#10 counter$count = 37319;
	#10 counter$count = 37320;
	#10 counter$count = 37321;
	#10 counter$count = 37322;
	#10 counter$count = 37323;
	#10 counter$count = 37324;
	#10 counter$count = 37325;
	#10 counter$count = 37326;
	#10 counter$count = 37327;
	#10 counter$count = 37328;
	#10 counter$count = 37329;
	#10 counter$count = 37330;
	#10 counter$count = 37331;
	#10 counter$count = 37332;
	#10 counter$count = 37333;
	#10 counter$count = 37334;
	#10 counter$count = 37335;
	#10 counter$count = 37336;
	#10 counter$count = 37337;
	#10 counter$count = 37338;
	#10 counter$count = 37339;
	#10 counter$count = 37340;
	#10 counter$count = 37341;
	#10 counter$count = 37342;
	#10 counter$count = 37343;
	#10 counter$count = 37344;
	#10 counter$count = 37345;
	#10 counter$count = 37346;
	#10 counter$count = 37347;
	#10 counter$count = 37348;
	#10 counter$count = 37349;
	#10 counter$count = 37350;
	#10 counter$count = 37351;
	#10 counter$count = 37352;
	#10 counter$count = 37353;
	#10 counter$count = 37354;
	#10 counter$count = 37355;
	#10 counter$count = 37356;
	#10 counter$count = 37357;
	#10 counter$count = 37358;
	#10 counter$count = 37359;
	#10 counter$count = 37360;
	#10 counter$count = 37361;
	#10 counter$count = 37362;
	#10 counter$count = 37363;
	#10 counter$count = 37364;
	#10 counter$count = 37365;
	#10 counter$count = 37366;
	#10 counter$count = 37367;
	#10 counter$count = 37368;
	#10 counter$count = 37369;
	#10 counter$count = 37370;
	#10 counter$count = 37371;
	#10 counter$count = 37372;
	#10 counter$count = 37373;
	#10 counter$count = 37374;
	#10 counter$count = 37375;
	#10 counter$count = 37376;
	#10 counter$count = 37377;
	#10 counter$count = 37378;
	#10 counter$count = 37379;
	#10 counter$count = 37380;
	#10 counter$count = 37381;
	#10 counter$count = 37382;
	#10 counter$count = 37383;
	#10 counter$count = 37384;
	#10 counter$count = 37385;
	#10 counter$count = 37386;
	#10 counter$count = 37387;
	#10 counter$count = 37388;
	#10 counter$count = 37389;
	#10 counter$count = 37390;
	#10 counter$count = 37391;
	#10 counter$count = 37392;
	#10 counter$count = 37393;
	#10 counter$count = 37394;
	#10 counter$count = 37395;
	#10 counter$count = 37396;
	#10 counter$count = 37397;
	#10 counter$count = 37398;
	#10 counter$count = 37399;
	#10 counter$count = 37400;
	#10 counter$count = 37401;
	#10 counter$count = 37402;
	#10 counter$count = 37403;
	#10 counter$count = 37404;
	#10 counter$count = 37405;
	#10 counter$count = 37406;
	#10 counter$count = 37407;
	#10 counter$count = 37408;
	#10 counter$count = 37409;
	#10 counter$count = 37410;
	#10 counter$count = 37411;
	#10 counter$count = 37412;
	#10 counter$count = 37413;
	#10 counter$count = 37414;
	#10 counter$count = 37415;
	#10 counter$count = 37416;
	#10 counter$count = 37417;
	#10 counter$count = 37418;
	#10 counter$count = 37419;
	#10 counter$count = 37420;
	#10 counter$count = 37421;
	#10 counter$count = 37422;
	#10 counter$count = 37423;
	#10 counter$count = 37424;
	#10 counter$count = 37425;
	#10 counter$count = 37426;
	#10 counter$count = 37427;
	#10 counter$count = 37428;
	#10 counter$count = 37429;
	#10 counter$count = 37430;
	#10 counter$count = 37431;
	#10 counter$count = 37432;
	#10 counter$count = 37433;
	#10 counter$count = 37434;
	#10 counter$count = 37435;
	#10 counter$count = 37436;
	#10 counter$count = 37437;
	#10 counter$count = 37438;
	#10 counter$count = 37439;
	#10 counter$count = 37440;
	#10 counter$count = 37441;
	#10 counter$count = 37442;
	#10 counter$count = 37443;
	#10 counter$count = 37444;
	#10 counter$count = 37445;
	#10 counter$count = 37446;
	#10 counter$count = 37447;
	#10 counter$count = 37448;
	#10 counter$count = 37449;
	#10 counter$count = 37450;
	#10 counter$count = 37451;
	#10 counter$count = 37452;
	#10 counter$count = 37453;
	#10 counter$count = 37454;
	#10 counter$count = 37455;
	#10 counter$count = 37456;
	#10 counter$count = 37457;
	#10 counter$count = 37458;
	#10 counter$count = 37459;
	#10 counter$count = 37460;
	#10 counter$count = 37461;
	#10 counter$count = 37462;
	#10 counter$count = 37463;
	#10 counter$count = 37464;
	#10 counter$count = 37465;
	#10 counter$count = 37466;
	#10 counter$count = 37467;
	#10 counter$count = 37468;
	#10 counter$count = 37469;
	#10 counter$count = 37470;
	#10 counter$count = 37471;
	#10 counter$count = 37472;
	#10 counter$count = 37473;
	#10 counter$count = 37474;
	#10 counter$count = 37475;
	#10 counter$count = 37476;
	#10 counter$count = 37477;
	#10 counter$count = 37478;
	#10 counter$count = 37479;
	#10 counter$count = 37480;
	#10 counter$count = 37481;
	#10 counter$count = 37482;
	#10 counter$count = 37483;
	#10 counter$count = 37484;
	#10 counter$count = 37485;
	#10 counter$count = 37486;
	#10 counter$count = 37487;
	#10 counter$count = 37488;
	#10 counter$count = 37489;
	#10 counter$count = 37490;
	#10 counter$count = 37491;
	#10 counter$count = 37492;
	#10 counter$count = 37493;
	#10 counter$count = 37494;
	#10 counter$count = 37495;
	#10 counter$count = 37496;
	#10 counter$count = 37497;
	#10 counter$count = 37498;
	#10 counter$count = 37499;
	#10 counter$count = 37500;
	#10 counter$count = 37501;
	#10 counter$count = 37502;
	#10 counter$count = 37503;
	#10 counter$count = 37504;
	#10 counter$count = 37505;
	#10 counter$count = 37506;
	#10 counter$count = 37507;
	#10 counter$count = 37508;
	#10 counter$count = 37509;
	#10 counter$count = 37510;
	#10 counter$count = 37511;
	#10 counter$count = 37512;
	#10 counter$count = 37513;
	#10 counter$count = 37514;
	#10 counter$count = 37515;
	#10 counter$count = 37516;
	#10 counter$count = 37517;
	#10 counter$count = 37518;
	#10 counter$count = 37519;
	#10 counter$count = 37520;
	#10 counter$count = 37521;
	#10 counter$count = 37522;
	#10 counter$count = 37523;
	#10 counter$count = 37524;
	#10 counter$count = 37525;
	#10 counter$count = 37526;
	#10 counter$count = 37527;
	#10 counter$count = 37528;
	#10 counter$count = 37529;
	#10 counter$count = 37530;
	#10 counter$count = 37531;
	#10 counter$count = 37532;
	#10 counter$count = 37533;
	#10 counter$count = 37534;
	#10 counter$count = 37535;
	#10 counter$count = 37536;
	#10 counter$count = 37537;
	#10 counter$count = 37538;
	#10 counter$count = 37539;
	#10 counter$count = 37540;
	#10 counter$count = 37541;
	#10 counter$count = 37542;
	#10 counter$count = 37543;
	#10 counter$count = 37544;
	#10 counter$count = 37545;
	#10 counter$count = 37546;
	#10 counter$count = 37547;
	#10 counter$count = 37548;
	#10 counter$count = 37549;
	#10 counter$count = 37550;
	#10 counter$count = 37551;
	#10 counter$count = 37552;
	#10 counter$count = 37553;
	#10 counter$count = 37554;
	#10 counter$count = 37555;
	#10 counter$count = 37556;
	#10 counter$count = 37557;
	#10 counter$count = 37558;
	#10 counter$count = 37559;
	#10 counter$count = 37560;
	#10 counter$count = 37561;
	#10 counter$count = 37562;
	#10 counter$count = 37563;
	#10 counter$count = 37564;
	#10 counter$count = 37565;
	#10 counter$count = 37566;
	#10 counter$count = 37567;
	#10 counter$count = 37568;
	#10 counter$count = 37569;
	#10 counter$count = 37570;
	#10 counter$count = 37571;
	#10 counter$count = 37572;
	#10 counter$count = 37573;
	#10 counter$count = 37574;
	#10 counter$count = 37575;
	#10 counter$count = 37576;
	#10 counter$count = 37577;
	#10 counter$count = 37578;
	#10 counter$count = 37579;
	#10 counter$count = 37580;
	#10 counter$count = 37581;
	#10 counter$count = 37582;
	#10 counter$count = 37583;
	#10 counter$count = 37584;
	#10 counter$count = 37585;
	#10 counter$count = 37586;
	#10 counter$count = 37587;
	#10 counter$count = 37588;
	#10 counter$count = 37589;
	#10 counter$count = 37590;
	#10 counter$count = 37591;
	#10 counter$count = 37592;
	#10 counter$count = 37593;
	#10 counter$count = 37594;
	#10 counter$count = 37595;
	#10 counter$count = 37596;
	#10 counter$count = 37597;
	#10 counter$count = 37598;
	#10 counter$count = 37599;
	#10 counter$count = 37600;
	#10 counter$count = 37601;
	#10 counter$count = 37602;
	#10 counter$count = 37603;
	#10 counter$count = 37604;
	#10 counter$count = 37605;
	#10 counter$count = 37606;
	#10 counter$count = 37607;
	#10 counter$count = 37608;
	#10 counter$count = 37609;
	#10 counter$count = 37610;
	#10 counter$count = 37611;
	#10 counter$count = 37612;
	#10 counter$count = 37613;
	#10 counter$count = 37614;
	#10 counter$count = 37615;
	#10 counter$count = 37616;
	#10 counter$count = 37617;
	#10 counter$count = 37618;
	#10 counter$count = 37619;
	#10 counter$count = 37620;
	#10 counter$count = 37621;
	#10 counter$count = 37622;
	#10 counter$count = 37623;
	#10 counter$count = 37624;
	#10 counter$count = 37625;
	#10 counter$count = 37626;
	#10 counter$count = 37627;
	#10 counter$count = 37628;
	#10 counter$count = 37629;
	#10 counter$count = 37630;
	#10 counter$count = 37631;
	#10 counter$count = 37632;
	#10 counter$count = 37633;
	#10 counter$count = 37634;
	#10 counter$count = 37635;
	#10 counter$count = 37636;
	#10 counter$count = 37637;
	#10 counter$count = 37638;
	#10 counter$count = 37639;
	#10 counter$count = 37640;
	#10 counter$count = 37641;
	#10 counter$count = 37642;
	#10 counter$count = 37643;
	#10 counter$count = 37644;
	#10 counter$count = 37645;
	#10 counter$count = 37646;
	#10 counter$count = 37647;
	#10 counter$count = 37648;
	#10 counter$count = 37649;
	#10 counter$count = 37650;
	#10 counter$count = 37651;
	#10 counter$count = 37652;
	#10 counter$count = 37653;
	#10 counter$count = 37654;
	#10 counter$count = 37655;
	#10 counter$count = 37656;
	#10 counter$count = 37657;
	#10 counter$count = 37658;
	#10 counter$count = 37659;
	#10 counter$count = 37660;
	#10 counter$count = 37661;
	#10 counter$count = 37662;
	#10 counter$count = 37663;
	#10 counter$count = 37664;
	#10 counter$count = 37665;
	#10 counter$count = 37666;
	#10 counter$count = 37667;
	#10 counter$count = 37668;
	#10 counter$count = 37669;
	#10 counter$count = 37670;
	#10 counter$count = 37671;
	#10 counter$count = 37672;
	#10 counter$count = 37673;
	#10 counter$count = 37674;
	#10 counter$count = 37675;
	#10 counter$count = 37676;
	#10 counter$count = 37677;
	#10 counter$count = 37678;
	#10 counter$count = 37679;
	#10 counter$count = 37680;
	#10 counter$count = 37681;
	#10 counter$count = 37682;
	#10 counter$count = 37683;
	#10 counter$count = 37684;
	#10 counter$count = 37685;
	#10 counter$count = 37686;
	#10 counter$count = 37687;
	#10 counter$count = 37688;
	#10 counter$count = 37689;
	#10 counter$count = 37690;
	#10 counter$count = 37691;
	#10 counter$count = 37692;
	#10 counter$count = 37693;
	#10 counter$count = 37694;
	#10 counter$count = 37695;
	#10 counter$count = 37696;
	#10 counter$count = 37697;
	#10 counter$count = 37698;
	#10 counter$count = 37699;
	#10 counter$count = 37700;
	#10 counter$count = 37701;
	#10 counter$count = 37702;
	#10 counter$count = 37703;
	#10 counter$count = 37704;
	#10 counter$count = 37705;
	#10 counter$count = 37706;
	#10 counter$count = 37707;
	#10 counter$count = 37708;
	#10 counter$count = 37709;
	#10 counter$count = 37710;
	#10 counter$count = 37711;
	#10 counter$count = 37712;
	#10 counter$count = 37713;
	#10 counter$count = 37714;
	#10 counter$count = 37715;
	#10 counter$count = 37716;
	#10 counter$count = 37717;
	#10 counter$count = 37718;
	#10 counter$count = 37719;
	#10 counter$count = 37720;
	#10 counter$count = 37721;
	#10 counter$count = 37722;
	#10 counter$count = 37723;
	#10 counter$count = 37724;
	#10 counter$count = 37725;
	#10 counter$count = 37726;
	#10 counter$count = 37727;
	#10 counter$count = 37728;
	#10 counter$count = 37729;
	#10 counter$count = 37730;
	#10 counter$count = 37731;
	#10 counter$count = 37732;
	#10 counter$count = 37733;
	#10 counter$count = 37734;
	#10 counter$count = 37735;
	#10 counter$count = 37736;
	#10 counter$count = 37737;
	#10 counter$count = 37738;
	#10 counter$count = 37739;
	#10 counter$count = 37740;
	#10 counter$count = 37741;
	#10 counter$count = 37742;
	#10 counter$count = 37743;
	#10 counter$count = 37744;
	#10 counter$count = 37745;
	#10 counter$count = 37746;
	#10 counter$count = 37747;
	#10 counter$count = 37748;
	#10 counter$count = 37749;
	#10 counter$count = 37750;
	#10 counter$count = 37751;
	#10 counter$count = 37752;
	#10 counter$count = 37753;
	#10 counter$count = 37754;
	#10 counter$count = 37755;
	#10 counter$count = 37756;
	#10 counter$count = 37757;
	#10 counter$count = 37758;
	#10 counter$count = 37759;
	#10 counter$count = 37760;
	#10 counter$count = 37761;
	#10 counter$count = 37762;
	#10 counter$count = 37763;
	#10 counter$count = 37764;
	#10 counter$count = 37765;
	#10 counter$count = 37766;
	#10 counter$count = 37767;
	#10 counter$count = 37768;
	#10 counter$count = 37769;
	#10 counter$count = 37770;
	#10 counter$count = 37771;
	#10 counter$count = 37772;
	#10 counter$count = 37773;
	#10 counter$count = 37774;
	#10 counter$count = 37775;
	#10 counter$count = 37776;
	#10 counter$count = 37777;
	#10 counter$count = 37778;
	#10 counter$count = 37779;
	#10 counter$count = 37780;
	#10 counter$count = 37781;
	#10 counter$count = 37782;
	#10 counter$count = 37783;
	#10 counter$count = 37784;
	#10 counter$count = 37785;
	#10 counter$count = 37786;
	#10 counter$count = 37787;
	#10 counter$count = 37788;
	#10 counter$count = 37789;
	#10 counter$count = 37790;
	#10 counter$count = 37791;
	#10 counter$count = 37792;
	#10 counter$count = 37793;
	#10 counter$count = 37794;
	#10 counter$count = 37795;
	#10 counter$count = 37796;
	#10 counter$count = 37797;
	#10 counter$count = 37798;
	#10 counter$count = 37799;
	#10 counter$count = 37800;
	#10 counter$count = 37801;
	#10 counter$count = 37802;
	#10 counter$count = 37803;
	#10 counter$count = 37804;
	#10 counter$count = 37805;
	#10 counter$count = 37806;
	#10 counter$count = 37807;
	#10 counter$count = 37808;
	#10 counter$count = 37809;
	#10 counter$count = 37810;
	#10 counter$count = 37811;
	#10 counter$count = 37812;
	#10 counter$count = 37813;
	#10 counter$count = 37814;
	#10 counter$count = 37815;
	#10 counter$count = 37816;
	#10 counter$count = 37817;
	#10 counter$count = 37818;
	#10 counter$count = 37819;
	#10 counter$count = 37820;
	#10 counter$count = 37821;
	#10 counter$count = 37822;
	#10 counter$count = 37823;
	#10 counter$count = 37824;
	#10 counter$count = 37825;
	#10 counter$count = 37826;
	#10 counter$count = 37827;
	#10 counter$count = 37828;
	#10 counter$count = 37829;
	#10 counter$count = 37830;
	#10 counter$count = 37831;
	#10 counter$count = 37832;
	#10 counter$count = 37833;
	#10 counter$count = 37834;
	#10 counter$count = 37835;
	#10 counter$count = 37836;
	#10 counter$count = 37837;
	#10 counter$count = 37838;
	#10 counter$count = 37839;
	#10 counter$count = 37840;
	#10 counter$count = 37841;
	#10 counter$count = 37842;
	#10 counter$count = 37843;
	#10 counter$count = 37844;
	#10 counter$count = 37845;
	#10 counter$count = 37846;
	#10 counter$count = 37847;
	#10 counter$count = 37848;
	#10 counter$count = 37849;
	#10 counter$count = 37850;
	#10 counter$count = 37851;
	#10 counter$count = 37852;
	#10 counter$count = 37853;
	#10 counter$count = 37854;
	#10 counter$count = 37855;
	#10 counter$count = 37856;
	#10 counter$count = 37857;
	#10 counter$count = 37858;
	#10 counter$count = 37859;
	#10 counter$count = 37860;
	#10 counter$count = 37861;
	#10 counter$count = 37862;
	#10 counter$count = 37863;
	#10 counter$count = 37864;
	#10 counter$count = 37865;
	#10 counter$count = 37866;
	#10 counter$count = 37867;
	#10 counter$count = 37868;
	#10 counter$count = 37869;
	#10 counter$count = 37870;
	#10 counter$count = 37871;
	#10 counter$count = 37872;
	#10 counter$count = 37873;
	#10 counter$count = 37874;
	#10 counter$count = 37875;
	#10 counter$count = 37876;
	#10 counter$count = 37877;
	#10 counter$count = 37878;
	#10 counter$count = 37879;
	#10 counter$count = 37880;
	#10 counter$count = 37881;
	#10 counter$count = 37882;
	#10 counter$count = 37883;
	#10 counter$count = 37884;
	#10 counter$count = 37885;
	#10 counter$count = 37886;
	#10 counter$count = 37887;
	#10 counter$count = 37888;
	#10 counter$count = 37889;
	#10 counter$count = 37890;
	#10 counter$count = 37891;
	#10 counter$count = 37892;
	#10 counter$count = 37893;
	#10 counter$count = 37894;
	#10 counter$count = 37895;
	#10 counter$count = 37896;
	#10 counter$count = 37897;
	#10 counter$count = 37898;
	#10 counter$count = 37899;
	#10 counter$count = 37900;
	#10 counter$count = 37901;
	#10 counter$count = 37902;
	#10 counter$count = 37903;
	#10 counter$count = 37904;
	#10 counter$count = 37905;
	#10 counter$count = 37906;
	#10 counter$count = 37907;
	#10 counter$count = 37908;
	#10 counter$count = 37909;
	#10 counter$count = 37910;
	#10 counter$count = 37911;
	#10 counter$count = 37912;
	#10 counter$count = 37913;
	#10 counter$count = 37914;
	#10 counter$count = 37915;
	#10 counter$count = 37916;
	#10 counter$count = 37917;
	#10 counter$count = 37918;
	#10 counter$count = 37919;
	#10 counter$count = 37920;
	#10 counter$count = 37921;
	#10 counter$count = 37922;
	#10 counter$count = 37923;
	#10 counter$count = 37924;
	#10 counter$count = 37925;
	#10 counter$count = 37926;
	#10 counter$count = 37927;
	#10 counter$count = 37928;
	#10 counter$count = 37929;
	#10 counter$count = 37930;
	#10 counter$count = 37931;
	#10 counter$count = 37932;
	#10 counter$count = 37933;
	#10 counter$count = 37934;
	#10 counter$count = 37935;
	#10 counter$count = 37936;
	#10 counter$count = 37937;
	#10 counter$count = 37938;
	#10 counter$count = 37939;
	#10 counter$count = 37940;
	#10 counter$count = 37941;
	#10 counter$count = 37942;
	#10 counter$count = 37943;
	#10 counter$count = 37944;
	#10 counter$count = 37945;
	#10 counter$count = 37946;
	#10 counter$count = 37947;
	#10 counter$count = 37948;
	#10 counter$count = 37949;
	#10 counter$count = 37950;
	#10 counter$count = 37951;
	#10 counter$count = 37952;
	#10 counter$count = 37953;
	#10 counter$count = 37954;
	#10 counter$count = 37955;
	#10 counter$count = 37956;
	#10 counter$count = 37957;
	#10 counter$count = 37958;
	#10 counter$count = 37959;
	#10 counter$count = 37960;
	#10 counter$count = 37961;
	#10 counter$count = 37962;
	#10 counter$count = 37963;
	#10 counter$count = 37964;
	#10 counter$count = 37965;
	#10 counter$count = 37966;
	#10 counter$count = 37967;
	#10 counter$count = 37968;
	#10 counter$count = 37969;
	#10 counter$count = 37970;
	#10 counter$count = 37971;
	#10 counter$count = 37972;
	#10 counter$count = 37973;
	#10 counter$count = 37974;
	#10 counter$count = 37975;
	#10 counter$count = 37976;
	#10 counter$count = 37977;
	#10 counter$count = 37978;
	#10 counter$count = 37979;
	#10 counter$count = 37980;
	#10 counter$count = 37981;
	#10 counter$count = 37982;
	#10 counter$count = 37983;
	#10 counter$count = 37984;
	#10 counter$count = 37985;
	#10 counter$count = 37986;
	#10 counter$count = 37987;
	#10 counter$count = 37988;
	#10 counter$count = 37989;
	#10 counter$count = 37990;
	#10 counter$count = 37991;
	#10 counter$count = 37992;
	#10 counter$count = 37993;
	#10 counter$count = 37994;
	#10 counter$count = 37995;
	#10 counter$count = 37996;
	#10 counter$count = 37997;
	#10 counter$count = 37998;
	#10 counter$count = 37999;
	#10 counter$count = 38000;
	#10 counter$count = 38001;
	#10 counter$count = 38002;
	#10 counter$count = 38003;
	#10 counter$count = 38004;
	#10 counter$count = 38005;
	#10 counter$count = 38006;
	#10 counter$count = 38007;
	#10 counter$count = 38008;
	#10 counter$count = 38009;
	#10 counter$count = 38010;
	#10 counter$count = 38011;
	#10 counter$count = 38012;
	#10 counter$count = 38013;
	#10 counter$count = 38014;
	#10 counter$count = 38015;
	#10 counter$count = 38016;
	#10 counter$count = 38017;
	#10 counter$count = 38018;
	#10 counter$count = 38019;
	#10 counter$count = 38020;
	#10 counter$count = 38021;
	#10 counter$count = 38022;
	#10 counter$count = 38023;
	#10 counter$count = 38024;
	#10 counter$count = 38025;
	#10 counter$count = 38026;
	#10 counter$count = 38027;
	#10 counter$count = 38028;
	#10 counter$count = 38029;
	#10 counter$count = 38030;
	#10 counter$count = 38031;
	#10 counter$count = 38032;
	#10 counter$count = 38033;
	#10 counter$count = 38034;
	#10 counter$count = 38035;
	#10 counter$count = 38036;
	#10 counter$count = 38037;
	#10 counter$count = 38038;
	#10 counter$count = 38039;
	#10 counter$count = 38040;
	#10 counter$count = 38041;
	#10 counter$count = 38042;
	#10 counter$count = 38043;
	#10 counter$count = 38044;
	#10 counter$count = 38045;
	#10 counter$count = 38046;
	#10 counter$count = 38047;
	#10 counter$count = 38048;
	#10 counter$count = 38049;
	#10 counter$count = 38050;
	#10 counter$count = 38051;
	#10 counter$count = 38052;
	#10 counter$count = 38053;
	#10 counter$count = 38054;
	#10 counter$count = 38055;
	#10 counter$count = 38056;
	#10 counter$count = 38057;
	#10 counter$count = 38058;
	#10 counter$count = 38059;
	#10 counter$count = 38060;
	#10 counter$count = 38061;
	#10 counter$count = 38062;
	#10 counter$count = 38063;
	#10 counter$count = 38064;
	#10 counter$count = 38065;
	#10 counter$count = 38066;
	#10 counter$count = 38067;
	#10 counter$count = 38068;
	#10 counter$count = 38069;
	#10 counter$count = 38070;
	#10 counter$count = 38071;
	#10 counter$count = 38072;
	#10 counter$count = 38073;
	#10 counter$count = 38074;
	#10 counter$count = 38075;
	#10 counter$count = 38076;
	#10 counter$count = 38077;
	#10 counter$count = 38078;
	#10 counter$count = 38079;
	#10 counter$count = 38080;
	#10 counter$count = 38081;
	#10 counter$count = 38082;
	#10 counter$count = 38083;
	#10 counter$count = 38084;
	#10 counter$count = 38085;
	#10 counter$count = 38086;
	#10 counter$count = 38087;
	#10 counter$count = 38088;
	#10 counter$count = 38089;
	#10 counter$count = 38090;
	#10 counter$count = 38091;
	#10 counter$count = 38092;
	#10 counter$count = 38093;
	#10 counter$count = 38094;
	#10 counter$count = 38095;
	#10 counter$count = 38096;
	#10 counter$count = 38097;
	#10 counter$count = 38098;
	#10 counter$count = 38099;
	#10 counter$count = 38100;
	#10 counter$count = 38101;
	#10 counter$count = 38102;
	#10 counter$count = 38103;
	#10 counter$count = 38104;
	#10 counter$count = 38105;
	#10 counter$count = 38106;
	#10 counter$count = 38107;
	#10 counter$count = 38108;
	#10 counter$count = 38109;
	#10 counter$count = 38110;
	#10 counter$count = 38111;
	#10 counter$count = 38112;
	#10 counter$count = 38113;
	#10 counter$count = 38114;
	#10 counter$count = 38115;
	#10 counter$count = 38116;
	#10 counter$count = 38117;
	#10 counter$count = 38118;
	#10 counter$count = 38119;
	#10 counter$count = 38120;
	#10 counter$count = 38121;
	#10 counter$count = 38122;
	#10 counter$count = 38123;
	#10 counter$count = 38124;
	#10 counter$count = 38125;
	#10 counter$count = 38126;
	#10 counter$count = 38127;
	#10 counter$count = 38128;
	#10 counter$count = 38129;
	#10 counter$count = 38130;
	#10 counter$count = 38131;
	#10 counter$count = 38132;
	#10 counter$count = 38133;
	#10 counter$count = 38134;
	#10 counter$count = 38135;
	#10 counter$count = 38136;
	#10 counter$count = 38137;
	#10 counter$count = 38138;
	#10 counter$count = 38139;
	#10 counter$count = 38140;
	#10 counter$count = 38141;
	#10 counter$count = 38142;
	#10 counter$count = 38143;
	#10 counter$count = 38144;
	#10 counter$count = 38145;
	#10 counter$count = 38146;
	#10 counter$count = 38147;
	#10 counter$count = 38148;
	#10 counter$count = 38149;
	#10 counter$count = 38150;
	#10 counter$count = 38151;
	#10 counter$count = 38152;
	#10 counter$count = 38153;
	#10 counter$count = 38154;
	#10 counter$count = 38155;
	#10 counter$count = 38156;
	#10 counter$count = 38157;
	#10 counter$count = 38158;
	#10 counter$count = 38159;
	#10 counter$count = 38160;
	#10 counter$count = 38161;
	#10 counter$count = 38162;
	#10 counter$count = 38163;
	#10 counter$count = 38164;
	#10 counter$count = 38165;
	#10 counter$count = 38166;
	#10 counter$count = 38167;
	#10 counter$count = 38168;
	#10 counter$count = 38169;
	#10 counter$count = 38170;
	#10 counter$count = 38171;
	#10 counter$count = 38172;
	#10 counter$count = 38173;
	#10 counter$count = 38174;
	#10 counter$count = 38175;
	#10 counter$count = 38176;
	#10 counter$count = 38177;
	#10 counter$count = 38178;
	#10 counter$count = 38179;
	#10 counter$count = 38180;
	#10 counter$count = 38181;
	#10 counter$count = 38182;
	#10 counter$count = 38183;
	#10 counter$count = 38184;
	#10 counter$count = 38185;
	#10 counter$count = 38186;
	#10 counter$count = 38187;
	#10 counter$count = 38188;
	#10 counter$count = 38189;
	#10 counter$count = 38190;
	#10 counter$count = 38191;
	#10 counter$count = 38192;
	#10 counter$count = 38193;
	#10 counter$count = 38194;
	#10 counter$count = 38195;
	#10 counter$count = 38196;
	#10 counter$count = 38197;
	#10 counter$count = 38198;
	#10 counter$count = 38199;
	#10 counter$count = 38200;
	#10 counter$count = 38201;
	#10 counter$count = 38202;
	#10 counter$count = 38203;
	#10 counter$count = 38204;
	#10 counter$count = 38205;
	#10 counter$count = 38206;
	#10 counter$count = 38207;
	#10 counter$count = 38208;
	#10 counter$count = 38209;
	#10 counter$count = 38210;
	#10 counter$count = 38211;
	#10 counter$count = 38212;
	#10 counter$count = 38213;
	#10 counter$count = 38214;
	#10 counter$count = 38215;
	#10 counter$count = 38216;
	#10 counter$count = 38217;
	#10 counter$count = 38218;
	#10 counter$count = 38219;
	#10 counter$count = 38220;
	#10 counter$count = 38221;
	#10 counter$count = 38222;
	#10 counter$count = 38223;
	#10 counter$count = 38224;
	#10 counter$count = 38225;
	#10 counter$count = 38226;
	#10 counter$count = 38227;
	#10 counter$count = 38228;
	#10 counter$count = 38229;
	#10 counter$count = 38230;
	#10 counter$count = 38231;
	#10 counter$count = 38232;
	#10 counter$count = 38233;
	#10 counter$count = 38234;
	#10 counter$count = 38235;
	#10 counter$count = 38236;
	#10 counter$count = 38237;
	#10 counter$count = 38238;
	#10 counter$count = 38239;
	#10 counter$count = 38240;
	#10 counter$count = 38241;
	#10 counter$count = 38242;
	#10 counter$count = 38243;
	#10 counter$count = 38244;
	#10 counter$count = 38245;
	#10 counter$count = 38246;
	#10 counter$count = 38247;
	#10 counter$count = 38248;
	#10 counter$count = 38249;
	#10 counter$count = 38250;
	#10 counter$count = 38251;
	#10 counter$count = 38252;
	#10 counter$count = 38253;
	#10 counter$count = 38254;
	#10 counter$count = 38255;
	#10 counter$count = 38256;
	#10 counter$count = 38257;
	#10 counter$count = 38258;
	#10 counter$count = 38259;
	#10 counter$count = 38260;
	#10 counter$count = 38261;
	#10 counter$count = 38262;
	#10 counter$count = 38263;
	#10 counter$count = 38264;
	#10 counter$count = 38265;
	#10 counter$count = 38266;
	#10 counter$count = 38267;
	#10 counter$count = 38268;
	#10 counter$count = 38269;
	#10 counter$count = 38270;
	#10 counter$count = 38271;
	#10 counter$count = 38272;
	#10 counter$count = 38273;
	#10 counter$count = 38274;
	#10 counter$count = 38275;
	#10 counter$count = 38276;
	#10 counter$count = 38277;
	#10 counter$count = 38278;
	#10 counter$count = 38279;
	#10 counter$count = 38280;
	#10 counter$count = 38281;
	#10 counter$count = 38282;
	#10 counter$count = 38283;
	#10 counter$count = 38284;
	#10 counter$count = 38285;
	#10 counter$count = 38286;
	#10 counter$count = 38287;
	#10 counter$count = 38288;
	#10 counter$count = 38289;
	#10 counter$count = 38290;
	#10 counter$count = 38291;
	#10 counter$count = 38292;
	#10 counter$count = 38293;
	#10 counter$count = 38294;
	#10 counter$count = 38295;
	#10 counter$count = 38296;
	#10 counter$count = 38297;
	#10 counter$count = 38298;
	#10 counter$count = 38299;
	#10 counter$count = 38300;
	#10 counter$count = 38301;
	#10 counter$count = 38302;
	#10 counter$count = 38303;
	#10 counter$count = 38304;
	#10 counter$count = 38305;
	#10 counter$count = 38306;
	#10 counter$count = 38307;
	#10 counter$count = 38308;
	#10 counter$count = 38309;
	#10 counter$count = 38310;
	#10 counter$count = 38311;
	#10 counter$count = 38312;
	#10 counter$count = 38313;
	#10 counter$count = 38314;
	#10 counter$count = 38315;
	#10 counter$count = 38316;
	#10 counter$count = 38317;
	#10 counter$count = 38318;
	#10 counter$count = 38319;
	#10 counter$count = 38320;
	#10 counter$count = 38321;
	#10 counter$count = 38322;
	#10 counter$count = 38323;
	#10 counter$count = 38324;
	#10 counter$count = 38325;
	#10 counter$count = 38326;
	#10 counter$count = 38327;
	#10 counter$count = 38328;
	#10 counter$count = 38329;
	#10 counter$count = 38330;
	#10 counter$count = 38331;
	#10 counter$count = 38332;
	#10 counter$count = 38333;
	#10 counter$count = 38334;
	#10 counter$count = 38335;
	#10 counter$count = 38336;
	#10 counter$count = 38337;
	#10 counter$count = 38338;
	#10 counter$count = 38339;
	#10 counter$count = 38340;
	#10 counter$count = 38341;
	#10 counter$count = 38342;
	#10 counter$count = 38343;
	#10 counter$count = 38344;
	#10 counter$count = 38345;
	#10 counter$count = 38346;
	#10 counter$count = 38347;
	#10 counter$count = 38348;
	#10 counter$count = 38349;
	#10 counter$count = 38350;
	#10 counter$count = 38351;
	#10 counter$count = 38352;
	#10 counter$count = 38353;
	#10 counter$count = 38354;
	#10 counter$count = 38355;
	#10 counter$count = 38356;
	#10 counter$count = 38357;
	#10 counter$count = 38358;
	#10 counter$count = 38359;
	#10 counter$count = 38360;
	#10 counter$count = 38361;
	#10 counter$count = 38362;
	#10 counter$count = 38363;
	#10 counter$count = 38364;
	#10 counter$count = 38365;
	#10 counter$count = 38366;
	#10 counter$count = 38367;
	#10 counter$count = 38368;
	#10 counter$count = 38369;
	#10 counter$count = 38370;
	#10 counter$count = 38371;
	#10 counter$count = 38372;
	#10 counter$count = 38373;
	#10 counter$count = 38374;
	#10 counter$count = 38375;
	#10 counter$count = 38376;
	#10 counter$count = 38377;
	#10 counter$count = 38378;
	#10 counter$count = 38379;
	#10 counter$count = 38380;
	#10 counter$count = 38381;
	#10 counter$count = 38382;
	#10 counter$count = 38383;
	#10 counter$count = 38384;
	#10 counter$count = 38385;
	#10 counter$count = 38386;
	#10 counter$count = 38387;
	#10 counter$count = 38388;
	#10 counter$count = 38389;
	#10 counter$count = 38390;
	#10 counter$count = 38391;
	#10 counter$count = 38392;
	#10 counter$count = 38393;
	#10 counter$count = 38394;
	#10 counter$count = 38395;
	#10 counter$count = 38396;
	#10 counter$count = 38397;
	#10 counter$count = 38398;
	#10 counter$count = 38399;
	#10 counter$count = 38400;
	#10 counter$count = 38401;
	#10 counter$count = 38402;
	#10 counter$count = 38403;
	#10 counter$count = 38404;
	#10 counter$count = 38405;
	#10 counter$count = 38406;
	#10 counter$count = 38407;
	#10 counter$count = 38408;
	#10 counter$count = 38409;
	#10 counter$count = 38410;
	#10 counter$count = 38411;
	#10 counter$count = 38412;
	#10 counter$count = 38413;
	#10 counter$count = 38414;
	#10 counter$count = 38415;
	#10 counter$count = 38416;
	#10 counter$count = 38417;
	#10 counter$count = 38418;
	#10 counter$count = 38419;
	#10 counter$count = 38420;
	#10 counter$count = 38421;
	#10 counter$count = 38422;
	#10 counter$count = 38423;
	#10 counter$count = 38424;
	#10 counter$count = 38425;
	#10 counter$count = 38426;
	#10 counter$count = 38427;
	#10 counter$count = 38428;
	#10 counter$count = 38429;
	#10 counter$count = 38430;
	#10 counter$count = 38431;
	#10 counter$count = 38432;
	#10 counter$count = 38433;
	#10 counter$count = 38434;
	#10 counter$count = 38435;
	#10 counter$count = 38436;
	#10 counter$count = 38437;
	#10 counter$count = 38438;
	#10 counter$count = 38439;
	#10 counter$count = 38440;
	#10 counter$count = 38441;
	#10 counter$count = 38442;
	#10 counter$count = 38443;
	#10 counter$count = 38444;
	#10 counter$count = 38445;
	#10 counter$count = 38446;
	#10 counter$count = 38447;
	#10 counter$count = 38448;
	#10 counter$count = 38449;
	#10 counter$count = 38450;
	#10 counter$count = 38451;
	#10 counter$count = 38452;
	#10 counter$count = 38453;
	#10 counter$count = 38454;
	#10 counter$count = 38455;
	#10 counter$count = 38456;
	#10 counter$count = 38457;
	#10 counter$count = 38458;
	#10 counter$count = 38459;
	#10 counter$count = 38460;
	#10 counter$count = 38461;
	#10 counter$count = 38462;
	#10 counter$count = 38463;
	#10 counter$count = 38464;
	#10 counter$count = 38465;
	#10 counter$count = 38466;
	#10 counter$count = 38467;
	#10 counter$count = 38468;
	#10 counter$count = 38469;
	#10 counter$count = 38470;
	#10 counter$count = 38471;
	#10 counter$count = 38472;
	#10 counter$count = 38473;
	#10 counter$count = 38474;
	#10 counter$count = 38475;
	#10 counter$count = 38476;
	#10 counter$count = 38477;
	#10 counter$count = 38478;
	#10 counter$count = 38479;
	#10 counter$count = 38480;
	#10 counter$count = 38481;
	#10 counter$count = 38482;
	#10 counter$count = 38483;
	#10 counter$count = 38484;
	#10 counter$count = 38485;
	#10 counter$count = 38486;
	#10 counter$count = 38487;
	#10 counter$count = 38488;
	#10 counter$count = 38489;
	#10 counter$count = 38490;
	#10 counter$count = 38491;
	#10 counter$count = 38492;
	#10 counter$count = 38493;
	#10 counter$count = 38494;
	#10 counter$count = 38495;
	#10 counter$count = 38496;
	#10 counter$count = 38497;
	#10 counter$count = 38498;
	#10 counter$count = 38499;
	#10 counter$count = 38500;
	#10 counter$count = 38501;
	#10 counter$count = 38502;
	#10 counter$count = 38503;
	#10 counter$count = 38504;
	#10 counter$count = 38505;
	#10 counter$count = 38506;
	#10 counter$count = 38507;
	#10 counter$count = 38508;
	#10 counter$count = 38509;
	#10 counter$count = 38510;
	#10 counter$count = 38511;
	#10 counter$count = 38512;
	#10 counter$count = 38513;
	#10 counter$count = 38514;
	#10 counter$count = 38515;
	#10 counter$count = 38516;
	#10 counter$count = 38517;
	#10 counter$count = 38518;
	#10 counter$count = 38519;
	#10 counter$count = 38520;
	#10 counter$count = 38521;
	#10 counter$count = 38522;
	#10 counter$count = 38523;
	#10 counter$count = 38524;
	#10 counter$count = 38525;
	#10 counter$count = 38526;
	#10 counter$count = 38527;
	#10 counter$count = 38528;
	#10 counter$count = 38529;
	#10 counter$count = 38530;
	#10 counter$count = 38531;
	#10 counter$count = 38532;
	#10 counter$count = 38533;
	#10 counter$count = 38534;
	#10 counter$count = 38535;
	#10 counter$count = 38536;
	#10 counter$count = 38537;
	#10 counter$count = 38538;
	#10 counter$count = 38539;
	#10 counter$count = 38540;
	#10 counter$count = 38541;
	#10 counter$count = 38542;
	#10 counter$count = 38543;
	#10 counter$count = 38544;
	#10 counter$count = 38545;
	#10 counter$count = 38546;
	#10 counter$count = 38547;
	#10 counter$count = 38548;
	#10 counter$count = 38549;
	#10 counter$count = 38550;
	#10 counter$count = 38551;
	#10 counter$count = 38552;
	#10 counter$count = 38553;
	#10 counter$count = 38554;
	#10 counter$count = 38555;
	#10 counter$count = 38556;
	#10 counter$count = 38557;
	#10 counter$count = 38558;
	#10 counter$count = 38559;
	#10 counter$count = 38560;
	#10 counter$count = 38561;
	#10 counter$count = 38562;
	#10 counter$count = 38563;
	#10 counter$count = 38564;
	#10 counter$count = 38565;
	#10 counter$count = 38566;
	#10 counter$count = 38567;
	#10 counter$count = 38568;
	#10 counter$count = 38569;
	#10 counter$count = 38570;
	#10 counter$count = 38571;
	#10 counter$count = 38572;
	#10 counter$count = 38573;
	#10 counter$count = 38574;
	#10 counter$count = 38575;
	#10 counter$count = 38576;
	#10 counter$count = 38577;
	#10 counter$count = 38578;
	#10 counter$count = 38579;
	#10 counter$count = 38580;
	#10 counter$count = 38581;
	#10 counter$count = 38582;
	#10 counter$count = 38583;
	#10 counter$count = 38584;
	#10 counter$count = 38585;
	#10 counter$count = 38586;
	#10 counter$count = 38587;
	#10 counter$count = 38588;
	#10 counter$count = 38589;
	#10 counter$count = 38590;
	#10 counter$count = 38591;
	#10 counter$count = 38592;
	#10 counter$count = 38593;
	#10 counter$count = 38594;
	#10 counter$count = 38595;
	#10 counter$count = 38596;
	#10 counter$count = 38597;
	#10 counter$count = 38598;
	#10 counter$count = 38599;
	#10 counter$count = 38600;
	#10 counter$count = 38601;
	#10 counter$count = 38602;
	#10 counter$count = 38603;
	#10 counter$count = 38604;
	#10 counter$count = 38605;
	#10 counter$count = 38606;
	#10 counter$count = 38607;
	#10 counter$count = 38608;
	#10 counter$count = 38609;
	#10 counter$count = 38610;
	#10 counter$count = 38611;
	#10 counter$count = 38612;
	#10 counter$count = 38613;
	#10 counter$count = 38614;
	#10 counter$count = 38615;
	#10 counter$count = 38616;
	#10 counter$count = 38617;
	#10 counter$count = 38618;
	#10 counter$count = 38619;
	#10 counter$count = 38620;
	#10 counter$count = 38621;
	#10 counter$count = 38622;
	#10 counter$count = 38623;
	#10 counter$count = 38624;
	#10 counter$count = 38625;
	#10 counter$count = 38626;
	#10 counter$count = 38627;
	#10 counter$count = 38628;
	#10 counter$count = 38629;
	#10 counter$count = 38630;
	#10 counter$count = 38631;
	#10 counter$count = 38632;
	#10 counter$count = 38633;
	#10 counter$count = 38634;
	#10 counter$count = 38635;
	#10 counter$count = 38636;
	#10 counter$count = 38637;
	#10 counter$count = 38638;
	#10 counter$count = 38639;
	#10 counter$count = 38640;
	#10 counter$count = 38641;
	#10 counter$count = 38642;
	#10 counter$count = 38643;
	#10 counter$count = 38644;
	#10 counter$count = 38645;
	#10 counter$count = 38646;
	#10 counter$count = 38647;
	#10 counter$count = 38648;
	#10 counter$count = 38649;
	#10 counter$count = 38650;
	#10 counter$count = 38651;
	#10 counter$count = 38652;
	#10 counter$count = 38653;
	#10 counter$count = 38654;
	#10 counter$count = 38655;
	#10 counter$count = 38656;
	#10 counter$count = 38657;
	#10 counter$count = 38658;
	#10 counter$count = 38659;
	#10 counter$count = 38660;
	#10 counter$count = 38661;
	#10 counter$count = 38662;
	#10 counter$count = 38663;
	#10 counter$count = 38664;
	#10 counter$count = 38665;
	#10 counter$count = 38666;
	#10 counter$count = 38667;
	#10 counter$count = 38668;
	#10 counter$count = 38669;
	#10 counter$count = 38670;
	#10 counter$count = 38671;
	#10 counter$count = 38672;
	#10 counter$count = 38673;
	#10 counter$count = 38674;
	#10 counter$count = 38675;
	#10 counter$count = 38676;
	#10 counter$count = 38677;
	#10 counter$count = 38678;
	#10 counter$count = 38679;
	#10 counter$count = 38680;
	#10 counter$count = 38681;
	#10 counter$count = 38682;
	#10 counter$count = 38683;
	#10 counter$count = 38684;
	#10 counter$count = 38685;
	#10 counter$count = 38686;
	#10 counter$count = 38687;
	#10 counter$count = 38688;
	#10 counter$count = 38689;
	#10 counter$count = 38690;
	#10 counter$count = 38691;
	#10 counter$count = 38692;
	#10 counter$count = 38693;
	#10 counter$count = 38694;
	#10 counter$count = 38695;
	#10 counter$count = 38696;
	#10 counter$count = 38697;
	#10 counter$count = 38698;
	#10 counter$count = 38699;
	#10 counter$count = 38700;
	#10 counter$count = 38701;
	#10 counter$count = 38702;
	#10 counter$count = 38703;
	#10 counter$count = 38704;
	#10 counter$count = 38705;
	#10 counter$count = 38706;
	#10 counter$count = 38707;
	#10 counter$count = 38708;
	#10 counter$count = 38709;
	#10 counter$count = 38710;
	#10 counter$count = 38711;
	#10 counter$count = 38712;
	#10 counter$count = 38713;
	#10 counter$count = 38714;
	#10 counter$count = 38715;
	#10 counter$count = 38716;
	#10 counter$count = 38717;
	#10 counter$count = 38718;
	#10 counter$count = 38719;
	#10 counter$count = 38720;
	#10 counter$count = 38721;
	#10 counter$count = 38722;
	#10 counter$count = 38723;
	#10 counter$count = 38724;
	#10 counter$count = 38725;
	#10 counter$count = 38726;
	#10 counter$count = 38727;
	#10 counter$count = 38728;
	#10 counter$count = 38729;
	#10 counter$count = 38730;
	#10 counter$count = 38731;
	#10 counter$count = 38732;
	#10 counter$count = 38733;
	#10 counter$count = 38734;
	#10 counter$count = 38735;
	#10 counter$count = 38736;
	#10 counter$count = 38737;
	#10 counter$count = 38738;
	#10 counter$count = 38739;
	#10 counter$count = 38740;
	#10 counter$count = 38741;
	#10 counter$count = 38742;
	#10 counter$count = 38743;
	#10 counter$count = 38744;
	#10 counter$count = 38745;
	#10 counter$count = 38746;
	#10 counter$count = 38747;
	#10 counter$count = 38748;
	#10 counter$count = 38749;
	#10 counter$count = 38750;
	#10 counter$count = 38751;
	#10 counter$count = 38752;
	#10 counter$count = 38753;
	#10 counter$count = 38754;
	#10 counter$count = 38755;
	#10 counter$count = 38756;
	#10 counter$count = 38757;
	#10 counter$count = 38758;
	#10 counter$count = 38759;
	#10 counter$count = 38760;
	#10 counter$count = 38761;
	#10 counter$count = 38762;
	#10 counter$count = 38763;
	#10 counter$count = 38764;
	#10 counter$count = 38765;
	#10 counter$count = 38766;
	#10 counter$count = 38767;
	#10 counter$count = 38768;
	#10 counter$count = 38769;
	#10 counter$count = 38770;
	#10 counter$count = 38771;
	#10 counter$count = 38772;
	#10 counter$count = 38773;
	#10 counter$count = 38774;
	#10 counter$count = 38775;
	#10 counter$count = 38776;
	#10 counter$count = 38777;
	#10 counter$count = 38778;
	#10 counter$count = 38779;
	#10 counter$count = 38780;
	#10 counter$count = 38781;
	#10 counter$count = 38782;
	#10 counter$count = 38783;
	#10 counter$count = 38784;
	#10 counter$count = 38785;
	#10 counter$count = 38786;
	#10 counter$count = 38787;
	#10 counter$count = 38788;
	#10 counter$count = 38789;
	#10 counter$count = 38790;
	#10 counter$count = 38791;
	#10 counter$count = 38792;
	#10 counter$count = 38793;
	#10 counter$count = 38794;
	#10 counter$count = 38795;
	#10 counter$count = 38796;
	#10 counter$count = 38797;
	#10 counter$count = 38798;
	#10 counter$count = 38799;
	#10 counter$count = 38800;
	#10 counter$count = 38801;
	#10 counter$count = 38802;
	#10 counter$count = 38803;
	#10 counter$count = 38804;
	#10 counter$count = 38805;
	#10 counter$count = 38806;
	#10 counter$count = 38807;
	#10 counter$count = 38808;
	#10 counter$count = 38809;
	#10 counter$count = 38810;
	#10 counter$count = 38811;
	#10 counter$count = 38812;
	#10 counter$count = 38813;
	#10 counter$count = 38814;
	#10 counter$count = 38815;
	#10 counter$count = 38816;
	#10 counter$count = 38817;
	#10 counter$count = 38818;
	#10 counter$count = 38819;
	#10 counter$count = 38820;
	#10 counter$count = 38821;
	#10 counter$count = 38822;
	#10 counter$count = 38823;
	#10 counter$count = 38824;
	#10 counter$count = 38825;
	#10 counter$count = 38826;
	#10 counter$count = 38827;
	#10 counter$count = 38828;
	#10 counter$count = 38829;
	#10 counter$count = 38830;
	#10 counter$count = 38831;
	#10 counter$count = 38832;
	#10 counter$count = 38833;
	#10 counter$count = 38834;
	#10 counter$count = 38835;
	#10 counter$count = 38836;
	#10 counter$count = 38837;
	#10 counter$count = 38838;
	#10 counter$count = 38839;
	#10 counter$count = 38840;
	#10 counter$count = 38841;
	#10 counter$count = 38842;
	#10 counter$count = 38843;
	#10 counter$count = 38844;
	#10 counter$count = 38845;
	#10 counter$count = 38846;
	#10 counter$count = 38847;
	#10 counter$count = 38848;
	#10 counter$count = 38849;
	#10 counter$count = 38850;
	#10 counter$count = 38851;
	#10 counter$count = 38852;
	#10 counter$count = 38853;
	#10 counter$count = 38854;
	#10 counter$count = 38855;
	#10 counter$count = 38856;
	#10 counter$count = 38857;
	#10 counter$count = 38858;
	#10 counter$count = 38859;
	#10 counter$count = 38860;
	#10 counter$count = 38861;
	#10 counter$count = 38862;
	#10 counter$count = 38863;
	#10 counter$count = 38864;
	#10 counter$count = 38865;
	#10 counter$count = 38866;
	#10 counter$count = 38867;
	#10 counter$count = 38868;
	#10 counter$count = 38869;
	#10 counter$count = 38870;
	#10 counter$count = 38871;
	#10 counter$count = 38872;
	#10 counter$count = 38873;
	#10 counter$count = 38874;
	#10 counter$count = 38875;
	#10 counter$count = 38876;
	#10 counter$count = 38877;
	#10 counter$count = 38878;
	#10 counter$count = 38879;
	#10 counter$count = 38880;
	#10 counter$count = 38881;
	#10 counter$count = 38882;
	#10 counter$count = 38883;
	#10 counter$count = 38884;
	#10 counter$count = 38885;
	#10 counter$count = 38886;
	#10 counter$count = 38887;
	#10 counter$count = 38888;
	#10 counter$count = 38889;
	#10 counter$count = 38890;
	#10 counter$count = 38891;
	#10 counter$count = 38892;
	#10 counter$count = 38893;
	#10 counter$count = 38894;
	#10 counter$count = 38895;
	#10 counter$count = 38896;
	#10 counter$count = 38897;
	#10 counter$count = 38898;
	#10 counter$count = 38899;
	#10 counter$count = 38900;
	#10 counter$count = 38901;
	#10 counter$count = 38902;
	#10 counter$count = 38903;
	#10 counter$count = 38904;
	#10 counter$count = 38905;
	#10 counter$count = 38906;
	#10 counter$count = 38907;
	#10 counter$count = 38908;
	#10 counter$count = 38909;
	#10 counter$count = 38910;
	#10 counter$count = 38911;
	#10 counter$count = 38912;
	#10 counter$count = 38913;
	#10 counter$count = 38914;
	#10 counter$count = 38915;
	#10 counter$count = 38916;
	#10 counter$count = 38917;
	#10 counter$count = 38918;
	#10 counter$count = 38919;
	#10 counter$count = 38920;
	#10 counter$count = 38921;
	#10 counter$count = 38922;
	#10 counter$count = 38923;
	#10 counter$count = 38924;
	#10 counter$count = 38925;
	#10 counter$count = 38926;
	#10 counter$count = 38927;
	#10 counter$count = 38928;
	#10 counter$count = 38929;
	#10 counter$count = 38930;
	#10 counter$count = 38931;
	#10 counter$count = 38932;
	#10 counter$count = 38933;
	#10 counter$count = 38934;
	#10 counter$count = 38935;
	#10 counter$count = 38936;
	#10 counter$count = 38937;
	#10 counter$count = 38938;
	#10 counter$count = 38939;
	#10 counter$count = 38940;
	#10 counter$count = 38941;
	#10 counter$count = 38942;
	#10 counter$count = 38943;
	#10 counter$count = 38944;
	#10 counter$count = 38945;
	#10 counter$count = 38946;
	#10 counter$count = 38947;
	#10 counter$count = 38948;
	#10 counter$count = 38949;
	#10 counter$count = 38950;
	#10 counter$count = 38951;
	#10 counter$count = 38952;
	#10 counter$count = 38953;
	#10 counter$count = 38954;
	#10 counter$count = 38955;
	#10 counter$count = 38956;
	#10 counter$count = 38957;
	#10 counter$count = 38958;
	#10 counter$count = 38959;
	#10 counter$count = 38960;
	#10 counter$count = 38961;
	#10 counter$count = 38962;
	#10 counter$count = 38963;
	#10 counter$count = 38964;
	#10 counter$count = 38965;
	#10 counter$count = 38966;
	#10 counter$count = 38967;
	#10 counter$count = 38968;
	#10 counter$count = 38969;
	#10 counter$count = 38970;
	#10 counter$count = 38971;
	#10 counter$count = 38972;
	#10 counter$count = 38973;
	#10 counter$count = 38974;
	#10 counter$count = 38975;
	#10 counter$count = 38976;
	#10 counter$count = 38977;
	#10 counter$count = 38978;
	#10 counter$count = 38979;
	#10 counter$count = 38980;
	#10 counter$count = 38981;
	#10 counter$count = 38982;
	#10 counter$count = 38983;
	#10 counter$count = 38984;
	#10 counter$count = 38985;
	#10 counter$count = 38986;
	#10 counter$count = 38987;
	#10 counter$count = 38988;
	#10 counter$count = 38989;
	#10 counter$count = 38990;
	#10 counter$count = 38991;
	#10 counter$count = 38992;
	#10 counter$count = 38993;
	#10 counter$count = 38994;
	#10 counter$count = 38995;
	#10 counter$count = 38996;
	#10 counter$count = 38997;
	#10 counter$count = 38998;
	#10 counter$count = 38999;
	#10 counter$count = 39000;
	#10 counter$count = 39001;
	#10 counter$count = 39002;
	#10 counter$count = 39003;
	#10 counter$count = 39004;
	#10 counter$count = 39005;
	#10 counter$count = 39006;
	#10 counter$count = 39007;
	#10 counter$count = 39008;
	#10 counter$count = 39009;
	#10 counter$count = 39010;
	#10 counter$count = 39011;
	#10 counter$count = 39012;
	#10 counter$count = 39013;
	#10 counter$count = 39014;
	#10 counter$count = 39015;
	#10 counter$count = 39016;
	#10 counter$count = 39017;
	#10 counter$count = 39018;
	#10 counter$count = 39019;
	#10 counter$count = 39020;
	#10 counter$count = 39021;
	#10 counter$count = 39022;
	#10 counter$count = 39023;
	#10 counter$count = 39024;
	#10 counter$count = 39025;
	#10 counter$count = 39026;
	#10 counter$count = 39027;
	#10 counter$count = 39028;
	#10 counter$count = 39029;
	#10 counter$count = 39030;
	#10 counter$count = 39031;
	#10 counter$count = 39032;
	#10 counter$count = 39033;
	#10 counter$count = 39034;
	#10 counter$count = 39035;
	#10 counter$count = 39036;
	#10 counter$count = 39037;
	#10 counter$count = 39038;
	#10 counter$count = 39039;
	#10 counter$count = 39040;
	#10 counter$count = 39041;
	#10 counter$count = 39042;
	#10 counter$count = 39043;
	#10 counter$count = 39044;
	#10 counter$count = 39045;
	#10 counter$count = 39046;
	#10 counter$count = 39047;
	#10 counter$count = 39048;
	#10 counter$count = 39049;
	#10 counter$count = 39050;
	#10 counter$count = 39051;
	#10 counter$count = 39052;
	#10 counter$count = 39053;
	#10 counter$count = 39054;
	#10 counter$count = 39055;
	#10 counter$count = 39056;
	#10 counter$count = 39057;
	#10 counter$count = 39058;
	#10 counter$count = 39059;
	#10 counter$count = 39060;
	#10 counter$count = 39061;
	#10 counter$count = 39062;
	#10 counter$count = 39063;
	#10 counter$count = 39064;
	#10 counter$count = 39065;
	#10 counter$count = 39066;
	#10 counter$count = 39067;
	#10 counter$count = 39068;
	#10 counter$count = 39069;
	#10 counter$count = 39070;
	#10 counter$count = 39071;
	#10 counter$count = 39072;
	#10 counter$count = 39073;
	#10 counter$count = 39074;
	#10 counter$count = 39075;
	#10 counter$count = 39076;
	#10 counter$count = 39077;
	#10 counter$count = 39078;
	#10 counter$count = 39079;
	#10 counter$count = 39080;
	#10 counter$count = 39081;
	#10 counter$count = 39082;
	#10 counter$count = 39083;
	#10 counter$count = 39084;
	#10 counter$count = 39085;
	#10 counter$count = 39086;
	#10 counter$count = 39087;
	#10 counter$count = 39088;
	#10 counter$count = 39089;
	#10 counter$count = 39090;
	#10 counter$count = 39091;
	#10 counter$count = 39092;
	#10 counter$count = 39093;
	#10 counter$count = 39094;
	#10 counter$count = 39095;
	#10 counter$count = 39096;
	#10 counter$count = 39097;
	#10 counter$count = 39098;
	#10 counter$count = 39099;
	#10 counter$count = 39100;
	#10 counter$count = 39101;
	#10 counter$count = 39102;
	#10 counter$count = 39103;
	#10 counter$count = 39104;
	#10 counter$count = 39105;
	#10 counter$count = 39106;
	#10 counter$count = 39107;
	#10 counter$count = 39108;
	#10 counter$count = 39109;
	#10 counter$count = 39110;
	#10 counter$count = 39111;
	#10 counter$count = 39112;
	#10 counter$count = 39113;
	#10 counter$count = 39114;
	#10 counter$count = 39115;
	#10 counter$count = 39116;
	#10 counter$count = 39117;
	#10 counter$count = 39118;
	#10 counter$count = 39119;
	#10 counter$count = 39120;
	#10 counter$count = 39121;
	#10 counter$count = 39122;
	#10 counter$count = 39123;
	#10 counter$count = 39124;
	#10 counter$count = 39125;
	#10 counter$count = 39126;
	#10 counter$count = 39127;
	#10 counter$count = 39128;
	#10 counter$count = 39129;
	#10 counter$count = 39130;
	#10 counter$count = 39131;
	#10 counter$count = 39132;
	#10 counter$count = 39133;
	#10 counter$count = 39134;
	#10 counter$count = 39135;
	#10 counter$count = 39136;
	#10 counter$count = 39137;
	#10 counter$count = 39138;
	#10 counter$count = 39139;
	#10 counter$count = 39140;
	#10 counter$count = 39141;
	#10 counter$count = 39142;
	#10 counter$count = 39143;
	#10 counter$count = 39144;
	#10 counter$count = 39145;
	#10 counter$count = 39146;
	#10 counter$count = 39147;
	#10 counter$count = 39148;
	#10 counter$count = 39149;
	#10 counter$count = 39150;
	#10 counter$count = 39151;
	#10 counter$count = 39152;
	#10 counter$count = 39153;
	#10 counter$count = 39154;
	#10 counter$count = 39155;
	#10 counter$count = 39156;
	#10 counter$count = 39157;
	#10 counter$count = 39158;
	#10 counter$count = 39159;
	#10 counter$count = 39160;
	#10 counter$count = 39161;
	#10 counter$count = 39162;
	#10 counter$count = 39163;
	#10 counter$count = 39164;
	#10 counter$count = 39165;
	#10 counter$count = 39166;
	#10 counter$count = 39167;
	#10 counter$count = 39168;
	#10 counter$count = 39169;
	#10 counter$count = 39170;
	#10 counter$count = 39171;
	#10 counter$count = 39172;
	#10 counter$count = 39173;
	#10 counter$count = 39174;
	#10 counter$count = 39175;
	#10 counter$count = 39176;
	#10 counter$count = 39177;
	#10 counter$count = 39178;
	#10 counter$count = 39179;
	#10 counter$count = 39180;
	#10 counter$count = 39181;
	#10 counter$count = 39182;
	#10 counter$count = 39183;
	#10 counter$count = 39184;
	#10 counter$count = 39185;
	#10 counter$count = 39186;
	#10 counter$count = 39187;
	#10 counter$count = 39188;
	#10 counter$count = 39189;
	#10 counter$count = 39190;
	#10 counter$count = 39191;
	#10 counter$count = 39192;
	#10 counter$count = 39193;
	#10 counter$count = 39194;
	#10 counter$count = 39195;
	#10 counter$count = 39196;
	#10 counter$count = 39197;
	#10 counter$count = 39198;
	#10 counter$count = 39199;
	#10 counter$count = 39200;
	#10 counter$count = 39201;
	#10 counter$count = 39202;
	#10 counter$count = 39203;
	#10 counter$count = 39204;
	#10 counter$count = 39205;
	#10 counter$count = 39206;
	#10 counter$count = 39207;
	#10 counter$count = 39208;
	#10 counter$count = 39209;
	#10 counter$count = 39210;
	#10 counter$count = 39211;
	#10 counter$count = 39212;
	#10 counter$count = 39213;
	#10 counter$count = 39214;
	#10 counter$count = 39215;
	#10 counter$count = 39216;
	#10 counter$count = 39217;
	#10 counter$count = 39218;
	#10 counter$count = 39219;
	#10 counter$count = 39220;
	#10 counter$count = 39221;
	#10 counter$count = 39222;
	#10 counter$count = 39223;
	#10 counter$count = 39224;
	#10 counter$count = 39225;
	#10 counter$count = 39226;
	#10 counter$count = 39227;
	#10 counter$count = 39228;
	#10 counter$count = 39229;
	#10 counter$count = 39230;
	#10 counter$count = 39231;
	#10 counter$count = 39232;
	#10 counter$count = 39233;
	#10 counter$count = 39234;
	#10 counter$count = 39235;
	#10 counter$count = 39236;
	#10 counter$count = 39237;
	#10 counter$count = 39238;
	#10 counter$count = 39239;
	#10 counter$count = 39240;
	#10 counter$count = 39241;
	#10 counter$count = 39242;
	#10 counter$count = 39243;
	#10 counter$count = 39244;
	#10 counter$count = 39245;
	#10 counter$count = 39246;
	#10 counter$count = 39247;
	#10 counter$count = 39248;
	#10 counter$count = 39249;
	#10 counter$count = 39250;
	#10 counter$count = 39251;
	#10 counter$count = 39252;
	#10 counter$count = 39253;
	#10 counter$count = 39254;
	#10 counter$count = 39255;
	#10 counter$count = 39256;
	#10 counter$count = 39257;
	#10 counter$count = 39258;
	#10 counter$count = 39259;
	#10 counter$count = 39260;
	#10 counter$count = 39261;
	#10 counter$count = 39262;
	#10 counter$count = 39263;
	#10 counter$count = 39264;
	#10 counter$count = 39265;
	#10 counter$count = 39266;
	#10 counter$count = 39267;
	#10 counter$count = 39268;
	#10 counter$count = 39269;
	#10 counter$count = 39270;
	#10 counter$count = 39271;
	#10 counter$count = 39272;
	#10 counter$count = 39273;
	#10 counter$count = 39274;
	#10 counter$count = 39275;
	#10 counter$count = 39276;
	#10 counter$count = 39277;
	#10 counter$count = 39278;
	#10 counter$count = 39279;
	#10 counter$count = 39280;
	#10 counter$count = 39281;
	#10 counter$count = 39282;
	#10 counter$count = 39283;
	#10 counter$count = 39284;
	#10 counter$count = 39285;
	#10 counter$count = 39286;
	#10 counter$count = 39287;
	#10 counter$count = 39288;
	#10 counter$count = 39289;
	#10 counter$count = 39290;
	#10 counter$count = 39291;
	#10 counter$count = 39292;
	#10 counter$count = 39293;
	#10 counter$count = 39294;
	#10 counter$count = 39295;
	#10 counter$count = 39296;
	#10 counter$count = 39297;
	#10 counter$count = 39298;
	#10 counter$count = 39299;
	#10 counter$count = 39300;
	#10 counter$count = 39301;
	#10 counter$count = 39302;
	#10 counter$count = 39303;
	#10 counter$count = 39304;
	#10 counter$count = 39305;
	#10 counter$count = 39306;
	#10 counter$count = 39307;
	#10 counter$count = 39308;
	#10 counter$count = 39309;
	#10 counter$count = 39310;
	#10 counter$count = 39311;
	#10 counter$count = 39312;
	#10 counter$count = 39313;
	#10 counter$count = 39314;
	#10 counter$count = 39315;
	#10 counter$count = 39316;
	#10 counter$count = 39317;
	#10 counter$count = 39318;
	#10 counter$count = 39319;
	#10 counter$count = 39320;
	#10 counter$count = 39321;
	#10 counter$count = 39322;
	#10 counter$count = 39323;
	#10 counter$count = 39324;
	#10 counter$count = 39325;
	#10 counter$count = 39326;
	#10 counter$count = 39327;
	#10 counter$count = 39328;
	#10 counter$count = 39329;
	#10 counter$count = 39330;
	#10 counter$count = 39331;
	#10 counter$count = 39332;
	#10 counter$count = 39333;
	#10 counter$count = 39334;
	#10 counter$count = 39335;
	#10 counter$count = 39336;
	#10 counter$count = 39337;
	#10 counter$count = 39338;
	#10 counter$count = 39339;
	#10 counter$count = 39340;
	#10 counter$count = 39341;
	#10 counter$count = 39342;
	#10 counter$count = 39343;
	#10 counter$count = 39344;
	#10 counter$count = 39345;
	#10 counter$count = 39346;
	#10 counter$count = 39347;
	#10 counter$count = 39348;
	#10 counter$count = 39349;
	#10 counter$count = 39350;
	#10 counter$count = 39351;
	#10 counter$count = 39352;
	#10 counter$count = 39353;
	#10 counter$count = 39354;
	#10 counter$count = 39355;
	#10 counter$count = 39356;
	#10 counter$count = 39357;
	#10 counter$count = 39358;
	#10 counter$count = 39359;
	#10 counter$count = 39360;
	#10 counter$count = 39361;
	#10 counter$count = 39362;
	#10 counter$count = 39363;
	#10 counter$count = 39364;
	#10 counter$count = 39365;
	#10 counter$count = 39366;
	#10 counter$count = 39367;
	#10 counter$count = 39368;
	#10 counter$count = 39369;
	#10 counter$count = 39370;
	#10 counter$count = 39371;
	#10 counter$count = 39372;
	#10 counter$count = 39373;
	#10 counter$count = 39374;
	#10 counter$count = 39375;
	#10 counter$count = 39376;
	#10 counter$count = 39377;
	#10 counter$count = 39378;
	#10 counter$count = 39379;
	#10 counter$count = 39380;
	#10 counter$count = 39381;
	#10 counter$count = 39382;
	#10 counter$count = 39383;
	#10 counter$count = 39384;
	#10 counter$count = 39385;
	#10 counter$count = 39386;
	#10 counter$count = 39387;
	#10 counter$count = 39388;
	#10 counter$count = 39389;
	#10 counter$count = 39390;
	#10 counter$count = 39391;
	#10 counter$count = 39392;
	#10 counter$count = 39393;
	#10 counter$count = 39394;
	#10 counter$count = 39395;
	#10 counter$count = 39396;
	#10 counter$count = 39397;
	#10 counter$count = 39398;
	#10 counter$count = 39399;
	#10 counter$count = 39400;
	#10 counter$count = 39401;
	#10 counter$count = 39402;
	#10 counter$count = 39403;
	#10 counter$count = 39404;
	#10 counter$count = 39405;
	#10 counter$count = 39406;
	#10 counter$count = 39407;
	#10 counter$count = 39408;
	#10 counter$count = 39409;
	#10 counter$count = 39410;
	#10 counter$count = 39411;
	#10 counter$count = 39412;
	#10 counter$count = 39413;
	#10 counter$count = 39414;
	#10 counter$count = 39415;
	#10 counter$count = 39416;
	#10 counter$count = 39417;
	#10 counter$count = 39418;
	#10 counter$count = 39419;
	#10 counter$count = 39420;
	#10 counter$count = 39421;
	#10 counter$count = 39422;
	#10 counter$count = 39423;
	#10 counter$count = 39424;
	#10 counter$count = 39425;
	#10 counter$count = 39426;
	#10 counter$count = 39427;
	#10 counter$count = 39428;
	#10 counter$count = 39429;
	#10 counter$count = 39430;
	#10 counter$count = 39431;
	#10 counter$count = 39432;
	#10 counter$count = 39433;
	#10 counter$count = 39434;
	#10 counter$count = 39435;
	#10 counter$count = 39436;
	#10 counter$count = 39437;
	#10 counter$count = 39438;
	#10 counter$count = 39439;
	#10 counter$count = 39440;
	#10 counter$count = 39441;
	#10 counter$count = 39442;
	#10 counter$count = 39443;
	#10 counter$count = 39444;
	#10 counter$count = 39445;
	#10 counter$count = 39446;
	#10 counter$count = 39447;
	#10 counter$count = 39448;
	#10 counter$count = 39449;
	#10 counter$count = 39450;
	#10 counter$count = 39451;
	#10 counter$count = 39452;
	#10 counter$count = 39453;
	#10 counter$count = 39454;
	#10 counter$count = 39455;
	#10 counter$count = 39456;
	#10 counter$count = 39457;
	#10 counter$count = 39458;
	#10 counter$count = 39459;
	#10 counter$count = 39460;
	#10 counter$count = 39461;
	#10 counter$count = 39462;
	#10 counter$count = 39463;
	#10 counter$count = 39464;
	#10 counter$count = 39465;
	#10 counter$count = 39466;
	#10 counter$count = 39467;
	#10 counter$count = 39468;
	#10 counter$count = 39469;
	#10 counter$count = 39470;
	#10 counter$count = 39471;
	#10 counter$count = 39472;
	#10 counter$count = 39473;
	#10 counter$count = 39474;
	#10 counter$count = 39475;
	#10 counter$count = 39476;
	#10 counter$count = 39477;
	#10 counter$count = 39478;
	#10 counter$count = 39479;
	#10 counter$count = 39480;
	#10 counter$count = 39481;
	#10 counter$count = 39482;
	#10 counter$count = 39483;
	#10 counter$count = 39484;
	#10 counter$count = 39485;
	#10 counter$count = 39486;
	#10 counter$count = 39487;
	#10 counter$count = 39488;
	#10 counter$count = 39489;
	#10 counter$count = 39490;
	#10 counter$count = 39491;
	#10 counter$count = 39492;
	#10 counter$count = 39493;
	#10 counter$count = 39494;
	#10 counter$count = 39495;
	#10 counter$count = 39496;
	#10 counter$count = 39497;
	#10 counter$count = 39498;
	#10 counter$count = 39499;
	#10 counter$count = 39500;
	#10 counter$count = 39501;
	#10 counter$count = 39502;
	#10 counter$count = 39503;
	#10 counter$count = 39504;
	#10 counter$count = 39505;
	#10 counter$count = 39506;
	#10 counter$count = 39507;
	#10 counter$count = 39508;
	#10 counter$count = 39509;
	#10 counter$count = 39510;
	#10 counter$count = 39511;
	#10 counter$count = 39512;
	#10 counter$count = 39513;
	#10 counter$count = 39514;
	#10 counter$count = 39515;
	#10 counter$count = 39516;
	#10 counter$count = 39517;
	#10 counter$count = 39518;
	#10 counter$count = 39519;
	#10 counter$count = 39520;
	#10 counter$count = 39521;
	#10 counter$count = 39522;
	#10 counter$count = 39523;
	#10 counter$count = 39524;
	#10 counter$count = 39525;
	#10 counter$count = 39526;
	#10 counter$count = 39527;
	#10 counter$count = 39528;
	#10 counter$count = 39529;
	#10 counter$count = 39530;
	#10 counter$count = 39531;
	#10 counter$count = 39532;
	#10 counter$count = 39533;
	#10 counter$count = 39534;
	#10 counter$count = 39535;
	#10 counter$count = 39536;
	#10 counter$count = 39537;
	#10 counter$count = 39538;
	#10 counter$count = 39539;
	#10 counter$count = 39540;
	#10 counter$count = 39541;
	#10 counter$count = 39542;
	#10 counter$count = 39543;
	#10 counter$count = 39544;
	#10 counter$count = 39545;
	#10 counter$count = 39546;
	#10 counter$count = 39547;
	#10 counter$count = 39548;
	#10 counter$count = 39549;
	#10 counter$count = 39550;
	#10 counter$count = 39551;
	#10 counter$count = 39552;
	#10 counter$count = 39553;
	#10 counter$count = 39554;
	#10 counter$count = 39555;
	#10 counter$count = 39556;
	#10 counter$count = 39557;
	#10 counter$count = 39558;
	#10 counter$count = 39559;
	#10 counter$count = 39560;
	#10 counter$count = 39561;
	#10 counter$count = 39562;
	#10 counter$count = 39563;
	#10 counter$count = 39564;
	#10 counter$count = 39565;
	#10 counter$count = 39566;
	#10 counter$count = 39567;
	#10 counter$count = 39568;
	#10 counter$count = 39569;
	#10 counter$count = 39570;
	#10 counter$count = 39571;
	#10 counter$count = 39572;
	#10 counter$count = 39573;
	#10 counter$count = 39574;
	#10 counter$count = 39575;
	#10 counter$count = 39576;
	#10 counter$count = 39577;
	#10 counter$count = 39578;
	#10 counter$count = 39579;
	#10 counter$count = 39580;
	#10 counter$count = 39581;
	#10 counter$count = 39582;
	#10 counter$count = 39583;
	#10 counter$count = 39584;
	#10 counter$count = 39585;
	#10 counter$count = 39586;
	#10 counter$count = 39587;
	#10 counter$count = 39588;
	#10 counter$count = 39589;
	#10 counter$count = 39590;
	#10 counter$count = 39591;
	#10 counter$count = 39592;
	#10 counter$count = 39593;
	#10 counter$count = 39594;
	#10 counter$count = 39595;
	#10 counter$count = 39596;
	#10 counter$count = 39597;
	#10 counter$count = 39598;
	#10 counter$count = 39599;
	#10 counter$count = 39600;
	#10 counter$count = 39601;
	#10 counter$count = 39602;
	#10 counter$count = 39603;
	#10 counter$count = 39604;
	#10 counter$count = 39605;
	#10 counter$count = 39606;
	#10 counter$count = 39607;
	#10 counter$count = 39608;
	#10 counter$count = 39609;
	#10 counter$count = 39610;
	#10 counter$count = 39611;
	#10 counter$count = 39612;
	#10 counter$count = 39613;
	#10 counter$count = 39614;
	#10 counter$count = 39615;
	#10 counter$count = 39616;
	#10 counter$count = 39617;
	#10 counter$count = 39618;
	#10 counter$count = 39619;
	#10 counter$count = 39620;
	#10 counter$count = 39621;
	#10 counter$count = 39622;
	#10 counter$count = 39623;
	#10 counter$count = 39624;
	#10 counter$count = 39625;
	#10 counter$count = 39626;
	#10 counter$count = 39627;
	#10 counter$count = 39628;
	#10 counter$count = 39629;
	#10 counter$count = 39630;
	#10 counter$count = 39631;
	#10 counter$count = 39632;
	#10 counter$count = 39633;
	#10 counter$count = 39634;
	#10 counter$count = 39635;
	#10 counter$count = 39636;
	#10 counter$count = 39637;
	#10 counter$count = 39638;
	#10 counter$count = 39639;
	#10 counter$count = 39640;
	#10 counter$count = 39641;
	#10 counter$count = 39642;
	#10 counter$count = 39643;
	#10 counter$count = 39644;
	#10 counter$count = 39645;
	#10 counter$count = 39646;
	#10 counter$count = 39647;
	#10 counter$count = 39648;
	#10 counter$count = 39649;
	#10 counter$count = 39650;
	#10 counter$count = 39651;
	#10 counter$count = 39652;
	#10 counter$count = 39653;
	#10 counter$count = 39654;
	#10 counter$count = 39655;
	#10 counter$count = 39656;
	#10 counter$count = 39657;
	#10 counter$count = 39658;
	#10 counter$count = 39659;
	#10 counter$count = 39660;
	#10 counter$count = 39661;
	#10 counter$count = 39662;
	#10 counter$count = 39663;
	#10 counter$count = 39664;
	#10 counter$count = 39665;
	#10 counter$count = 39666;
	#10 counter$count = 39667;
	#10 counter$count = 39668;
	#10 counter$count = 39669;
	#10 counter$count = 39670;
	#10 counter$count = 39671;
	#10 counter$count = 39672;
	#10 counter$count = 39673;
	#10 counter$count = 39674;
	#10 counter$count = 39675;
	#10 counter$count = 39676;
	#10 counter$count = 39677;
	#10 counter$count = 39678;
	#10 counter$count = 39679;
	#10 counter$count = 39680;
	#10 counter$count = 39681;
	#10 counter$count = 39682;
	#10 counter$count = 39683;
	#10 counter$count = 39684;
	#10 counter$count = 39685;
	#10 counter$count = 39686;
	#10 counter$count = 39687;
	#10 counter$count = 39688;
	#10 counter$count = 39689;
	#10 counter$count = 39690;
	#10 counter$count = 39691;
	#10 counter$count = 39692;
	#10 counter$count = 39693;
	#10 counter$count = 39694;
	#10 counter$count = 39695;
	#10 counter$count = 39696;
	#10 counter$count = 39697;
	#10 counter$count = 39698;
	#10 counter$count = 39699;
	#10 counter$count = 39700;
	#10 counter$count = 39701;
	#10 counter$count = 39702;
	#10 counter$count = 39703;
	#10 counter$count = 39704;
	#10 counter$count = 39705;
	#10 counter$count = 39706;
	#10 counter$count = 39707;
	#10 counter$count = 39708;
	#10 counter$count = 39709;
	#10 counter$count = 39710;
	#10 counter$count = 39711;
	#10 counter$count = 39712;
	#10 counter$count = 39713;
	#10 counter$count = 39714;
	#10 counter$count = 39715;
	#10 counter$count = 39716;
	#10 counter$count = 39717;
	#10 counter$count = 39718;
	#10 counter$count = 39719;
	#10 counter$count = 39720;
	#10 counter$count = 39721;
	#10 counter$count = 39722;
	#10 counter$count = 39723;
	#10 counter$count = 39724;
	#10 counter$count = 39725;
	#10 counter$count = 39726;
	#10 counter$count = 39727;
	#10 counter$count = 39728;
	#10 counter$count = 39729;
	#10 counter$count = 39730;
	#10 counter$count = 39731;
	#10 counter$count = 39732;
	#10 counter$count = 39733;
	#10 counter$count = 39734;
	#10 counter$count = 39735;
	#10 counter$count = 39736;
	#10 counter$count = 39737;
	#10 counter$count = 39738;
	#10 counter$count = 39739;
	#10 counter$count = 39740;
	#10 counter$count = 39741;
	#10 counter$count = 39742;
	#10 counter$count = 39743;
	#10 counter$count = 39744;
	#10 counter$count = 39745;
	#10 counter$count = 39746;
	#10 counter$count = 39747;
	#10 counter$count = 39748;
	#10 counter$count = 39749;
	#10 counter$count = 39750;
	#10 counter$count = 39751;
	#10 counter$count = 39752;
	#10 counter$count = 39753;
	#10 counter$count = 39754;
	#10 counter$count = 39755;
	#10 counter$count = 39756;
	#10 counter$count = 39757;
	#10 counter$count = 39758;
	#10 counter$count = 39759;
	#10 counter$count = 39760;
	#10 counter$count = 39761;
	#10 counter$count = 39762;
	#10 counter$count = 39763;
	#10 counter$count = 39764;
	#10 counter$count = 39765;
	#10 counter$count = 39766;
	#10 counter$count = 39767;
	#10 counter$count = 39768;
	#10 counter$count = 39769;
	#10 counter$count = 39770;
	#10 counter$count = 39771;
	#10 counter$count = 39772;
	#10 counter$count = 39773;
	#10 counter$count = 39774;
	#10 counter$count = 39775;
	#10 counter$count = 39776;
	#10 counter$count = 39777;
	#10 counter$count = 39778;
	#10 counter$count = 39779;
	#10 counter$count = 39780;
	#10 counter$count = 39781;
	#10 counter$count = 39782;
	#10 counter$count = 39783;
	#10 counter$count = 39784;
	#10 counter$count = 39785;
	#10 counter$count = 39786;
	#10 counter$count = 39787;
	#10 counter$count = 39788;
	#10 counter$count = 39789;
	#10 counter$count = 39790;
	#10 counter$count = 39791;
	#10 counter$count = 39792;
	#10 counter$count = 39793;
	#10 counter$count = 39794;
	#10 counter$count = 39795;
	#10 counter$count = 39796;
	#10 counter$count = 39797;
	#10 counter$count = 39798;
	#10 counter$count = 39799;
	#10 counter$count = 39800;
	#10 counter$count = 39801;
	#10 counter$count = 39802;
	#10 counter$count = 39803;
	#10 counter$count = 39804;
	#10 counter$count = 39805;
	#10 counter$count = 39806;
	#10 counter$count = 39807;
	#10 counter$count = 39808;
	#10 counter$count = 39809;
	#10 counter$count = 39810;
	#10 counter$count = 39811;
	#10 counter$count = 39812;
	#10 counter$count = 39813;
	#10 counter$count = 39814;
	#10 counter$count = 39815;
	#10 counter$count = 39816;
	#10 counter$count = 39817;
	#10 counter$count = 39818;
	#10 counter$count = 39819;
	#10 counter$count = 39820;
	#10 counter$count = 39821;
	#10 counter$count = 39822;
	#10 counter$count = 39823;
	#10 counter$count = 39824;
	#10 counter$count = 39825;
	#10 counter$count = 39826;
	#10 counter$count = 39827;
	#10 counter$count = 39828;
	#10 counter$count = 39829;
	#10 counter$count = 39830;
	#10 counter$count = 39831;
	#10 counter$count = 39832;
	#10 counter$count = 39833;
	#10 counter$count = 39834;
	#10 counter$count = 39835;
	#10 counter$count = 39836;
	#10 counter$count = 39837;
	#10 counter$count = 39838;
	#10 counter$count = 39839;
	#10 counter$count = 39840;
	#10 counter$count = 39841;
	#10 counter$count = 39842;
	#10 counter$count = 39843;
	#10 counter$count = 39844;
	#10 counter$count = 39845;
	#10 counter$count = 39846;
	#10 counter$count = 39847;
	#10 counter$count = 39848;
	#10 counter$count = 39849;
	#10 counter$count = 39850;
	#10 counter$count = 39851;
	#10 counter$count = 39852;
	#10 counter$count = 39853;
	#10 counter$count = 39854;
	#10 counter$count = 39855;
	#10 counter$count = 39856;
	#10 counter$count = 39857;
	#10 counter$count = 39858;
	#10 counter$count = 39859;
	#10 counter$count = 39860;
	#10 counter$count = 39861;
	#10 counter$count = 39862;
	#10 counter$count = 39863;
	#10 counter$count = 39864;
	#10 counter$count = 39865;
	#10 counter$count = 39866;
	#10 counter$count = 39867;
	#10 counter$count = 39868;
	#10 counter$count = 39869;
	#10 counter$count = 39870;
	#10 counter$count = 39871;
	#10 counter$count = 39872;
	#10 counter$count = 39873;
	#10 counter$count = 39874;
	#10 counter$count = 39875;
	#10 counter$count = 39876;
	#10 counter$count = 39877;
	#10 counter$count = 39878;
	#10 counter$count = 39879;
	#10 counter$count = 39880;
	#10 counter$count = 39881;
	#10 counter$count = 39882;
	#10 counter$count = 39883;
	#10 counter$count = 39884;
	#10 counter$count = 39885;
	#10 counter$count = 39886;
	#10 counter$count = 39887;
	#10 counter$count = 39888;
	#10 counter$count = 39889;
	#10 counter$count = 39890;
	#10 counter$count = 39891;
	#10 counter$count = 39892;
	#10 counter$count = 39893;
	#10 counter$count = 39894;
	#10 counter$count = 39895;
	#10 counter$count = 39896;
	#10 counter$count = 39897;
	#10 counter$count = 39898;
	#10 counter$count = 39899;
	#10 counter$count = 39900;
	#10 counter$count = 39901;
	#10 counter$count = 39902;
	#10 counter$count = 39903;
	#10 counter$count = 39904;
	#10 counter$count = 39905;
	#10 counter$count = 39906;
	#10 counter$count = 39907;
	#10 counter$count = 39908;
	#10 counter$count = 39909;
	#10 counter$count = 39910;
	#10 counter$count = 39911;
	#10 counter$count = 39912;
	#10 counter$count = 39913;
	#10 counter$count = 39914;
	#10 counter$count = 39915;
	#10 counter$count = 39916;
	#10 counter$count = 39917;
	#10 counter$count = 39918;
	#10 counter$count = 39919;
	#10 counter$count = 39920;
	#10 counter$count = 39921;
	#10 counter$count = 39922;
	#10 counter$count = 39923;
	#10 counter$count = 39924;
	#10 counter$count = 39925;
	#10 counter$count = 39926;
	#10 counter$count = 39927;
	#10 counter$count = 39928;
	#10 counter$count = 39929;
	#10 counter$count = 39930;
	#10 counter$count = 39931;
	#10 counter$count = 39932;
	#10 counter$count = 39933;
	#10 counter$count = 39934;
	#10 counter$count = 39935;
	#10 counter$count = 39936;
	#10 counter$count = 39937;
	#10 counter$count = 39938;
	#10 counter$count = 39939;
	#10 counter$count = 39940;
	#10 counter$count = 39941;
	#10 counter$count = 39942;
	#10 counter$count = 39943;
	#10 counter$count = 39944;
	#10 counter$count = 39945;
	#10 counter$count = 39946;
	#10 counter$count = 39947;
	#10 counter$count = 39948;
	#10 counter$count = 39949;
	#10 counter$count = 39950;
	#10 counter$count = 39951;
	#10 counter$count = 39952;
	#10 counter$count = 39953;
	#10 counter$count = 39954;
	#10 counter$count = 39955;
	#10 counter$count = 39956;
	#10 counter$count = 39957;
	#10 counter$count = 39958;
	#10 counter$count = 39959;
	#10 counter$count = 39960;
	#10 counter$count = 39961;
	#10 counter$count = 39962;
	#10 counter$count = 39963;
	#10 counter$count = 39964;
	#10 counter$count = 39965;
	#10 counter$count = 39966;
	#10 counter$count = 39967;
	#10 counter$count = 39968;
	#10 counter$count = 39969;
	#10 counter$count = 39970;
	#10 counter$count = 39971;
	#10 counter$count = 39972;
	#10 counter$count = 39973;
	#10 counter$count = 39974;
	#10 counter$count = 39975;
	#10 counter$count = 39976;
	#10 counter$count = 39977;
	#10 counter$count = 39978;
	#10 counter$count = 39979;
	#10 counter$count = 39980;
	#10 counter$count = 39981;
	#10 counter$count = 39982;
	#10 counter$count = 39983;
	#10 counter$count = 39984;
	#10 counter$count = 39985;
	#10 counter$count = 39986;
	#10 counter$count = 39987;
	#10 counter$count = 39988;
	#10 counter$count = 39989;
	#10 counter$count = 39990;
	#10 counter$count = 39991;
	#10 counter$count = 39992;
	#10 counter$count = 39993;
	#10 counter$count = 39994;
	#10 counter$count = 39995;
	#10 counter$count = 39996;
	#10 counter$count = 39997;
	#10 counter$count = 39998;
	#10 counter$count = 39999;
	#10 counter$count = 40000;
	#10 counter$count = 40001;
	#10 counter$count = 40002;
	#10 counter$count = 40003;
	#10 counter$count = 40004;
	#10 counter$count = 40005;
	#10 counter$count = 40006;
	#10 counter$count = 40007;
	#10 counter$count = 40008;
	#10 counter$count = 40009;
	#10 counter$count = 40010;
	#10 counter$count = 40011;
	#10 counter$count = 40012;
	#10 counter$count = 40013;
	#10 counter$count = 40014;
	#10 counter$count = 40015;
	#10 counter$count = 40016;
	#10 counter$count = 40017;
	#10 counter$count = 40018;
	#10 counter$count = 40019;
	#10 counter$count = 40020;
	#10 counter$count = 40021;
	#10 counter$count = 40022;
	#10 counter$count = 40023;
	#10 counter$count = 40024;
	#10 counter$count = 40025;
	#10 counter$count = 40026;
	#10 counter$count = 40027;
	#10 counter$count = 40028;
	#10 counter$count = 40029;
	#10 counter$count = 40030;
	#10 counter$count = 40031;
	#10 counter$count = 40032;
	#10 counter$count = 40033;
	#10 counter$count = 40034;
	#10 counter$count = 40035;
	#10 counter$count = 40036;
	#10 counter$count = 40037;
	#10 counter$count = 40038;
	#10 counter$count = 40039;
	#10 counter$count = 40040;
	#10 counter$count = 40041;
	#10 counter$count = 40042;
	#10 counter$count = 40043;
	#10 counter$count = 40044;
	#10 counter$count = 40045;
	#10 counter$count = 40046;
	#10 counter$count = 40047;
	#10 counter$count = 40048;
	#10 counter$count = 40049;
	#10 counter$count = 40050;
	#10 counter$count = 40051;
	#10 counter$count = 40052;
	#10 counter$count = 40053;
	#10 counter$count = 40054;
	#10 counter$count = 40055;
	#10 counter$count = 40056;
	#10 counter$count = 40057;
	#10 counter$count = 40058;
	#10 counter$count = 40059;
	#10 counter$count = 40060;
	#10 counter$count = 40061;
	#10 counter$count = 40062;
	#10 counter$count = 40063;
	#10 counter$count = 40064;
	#10 counter$count = 40065;
	#10 counter$count = 40066;
	#10 counter$count = 40067;
	#10 counter$count = 40068;
	#10 counter$count = 40069;
	#10 counter$count = 40070;
	#10 counter$count = 40071;
	#10 counter$count = 40072;
	#10 counter$count = 40073;
	#10 counter$count = 40074;
	#10 counter$count = 40075;
	#10 counter$count = 40076;
	#10 counter$count = 40077;
	#10 counter$count = 40078;
	#10 counter$count = 40079;
	#10 counter$count = 40080;
	#10 counter$count = 40081;
	#10 counter$count = 40082;
	#10 counter$count = 40083;
	#10 counter$count = 40084;
	#10 counter$count = 40085;
	#10 counter$count = 40086;
	#10 counter$count = 40087;
	#10 counter$count = 40088;
	#10 counter$count = 40089;
	#10 counter$count = 40090;
	#10 counter$count = 40091;
	#10 counter$count = 40092;
	#10 counter$count = 40093;
	#10 counter$count = 40094;
	#10 counter$count = 40095;
	#10 counter$count = 40096;
	#10 counter$count = 40097;
	#10 counter$count = 40098;
	#10 counter$count = 40099;
	#10 counter$count = 40100;
	#10 counter$count = 40101;
	#10 counter$count = 40102;
	#10 counter$count = 40103;
	#10 counter$count = 40104;
	#10 counter$count = 40105;
	#10 counter$count = 40106;
	#10 counter$count = 40107;
	#10 counter$count = 40108;
	#10 counter$count = 40109;
	#10 counter$count = 40110;
	#10 counter$count = 40111;
	#10 counter$count = 40112;
	#10 counter$count = 40113;
	#10 counter$count = 40114;
	#10 counter$count = 40115;
	#10 counter$count = 40116;
	#10 counter$count = 40117;
	#10 counter$count = 40118;
	#10 counter$count = 40119;
	#10 counter$count = 40120;
	#10 counter$count = 40121;
	#10 counter$count = 40122;
	#10 counter$count = 40123;
	#10 counter$count = 40124;
	#10 counter$count = 40125;
	#10 counter$count = 40126;
	#10 counter$count = 40127;
	#10 counter$count = 40128;
	#10 counter$count = 40129;
	#10 counter$count = 40130;
	#10 counter$count = 40131;
	#10 counter$count = 40132;
	#10 counter$count = 40133;
	#10 counter$count = 40134;
	#10 counter$count = 40135;
	#10 counter$count = 40136;
	#10 counter$count = 40137;
	#10 counter$count = 40138;
	#10 counter$count = 40139;
	#10 counter$count = 40140;
	#10 counter$count = 40141;
	#10 counter$count = 40142;
	#10 counter$count = 40143;
	#10 counter$count = 40144;
	#10 counter$count = 40145;
	#10 counter$count = 40146;
	#10 counter$count = 40147;
	#10 counter$count = 40148;
	#10 counter$count = 40149;
	#10 counter$count = 40150;
	#10 counter$count = 40151;
	#10 counter$count = 40152;
	#10 counter$count = 40153;
	#10 counter$count = 40154;
	#10 counter$count = 40155;
	#10 counter$count = 40156;
	#10 counter$count = 40157;
	#10 counter$count = 40158;
	#10 counter$count = 40159;
	#10 counter$count = 40160;
	#10 counter$count = 40161;
	#10 counter$count = 40162;
	#10 counter$count = 40163;
	#10 counter$count = 40164;
	#10 counter$count = 40165;
	#10 counter$count = 40166;
	#10 counter$count = 40167;
	#10 counter$count = 40168;
	#10 counter$count = 40169;
	#10 counter$count = 40170;
	#10 counter$count = 40171;
	#10 counter$count = 40172;
	#10 counter$count = 40173;
	#10 counter$count = 40174;
	#10 counter$count = 40175;
	#10 counter$count = 40176;
	#10 counter$count = 40177;
	#10 counter$count = 40178;
	#10 counter$count = 40179;
	#10 counter$count = 40180;
	#10 counter$count = 40181;
	#10 counter$count = 40182;
	#10 counter$count = 40183;
	#10 counter$count = 40184;
	#10 counter$count = 40185;
	#10 counter$count = 40186;
	#10 counter$count = 40187;
	#10 counter$count = 40188;
	#10 counter$count = 40189;
	#10 counter$count = 40190;
	#10 counter$count = 40191;
	#10 counter$count = 40192;
	#10 counter$count = 40193;
	#10 counter$count = 40194;
	#10 counter$count = 40195;
	#10 counter$count = 40196;
	#10 counter$count = 40197;
	#10 counter$count = 40198;
	#10 counter$count = 40199;
	#10 counter$count = 40200;
	#10 counter$count = 40201;
	#10 counter$count = 40202;
	#10 counter$count = 40203;
	#10 counter$count = 40204;
	#10 counter$count = 40205;
	#10 counter$count = 40206;
	#10 counter$count = 40207;
	#10 counter$count = 40208;
	#10 counter$count = 40209;
	#10 counter$count = 40210;
	#10 counter$count = 40211;
	#10 counter$count = 40212;
	#10 counter$count = 40213;
	#10 counter$count = 40214;
	#10 counter$count = 40215;
	#10 counter$count = 40216;
	#10 counter$count = 40217;
	#10 counter$count = 40218;
	#10 counter$count = 40219;
	#10 counter$count = 40220;
	#10 counter$count = 40221;
	#10 counter$count = 40222;
	#10 counter$count = 40223;
	#10 counter$count = 40224;
	#10 counter$count = 40225;
	#10 counter$count = 40226;
	#10 counter$count = 40227;
	#10 counter$count = 40228;
	#10 counter$count = 40229;
	#10 counter$count = 40230;
	#10 counter$count = 40231;
	#10 counter$count = 40232;
	#10 counter$count = 40233;
	#10 counter$count = 40234;
	#10 counter$count = 40235;
	#10 counter$count = 40236;
	#10 counter$count = 40237;
	#10 counter$count = 40238;
	#10 counter$count = 40239;
	#10 counter$count = 40240;
	#10 counter$count = 40241;
	#10 counter$count = 40242;
	#10 counter$count = 40243;
	#10 counter$count = 40244;
	#10 counter$count = 40245;
	#10 counter$count = 40246;
	#10 counter$count = 40247;
	#10 counter$count = 40248;
	#10 counter$count = 40249;
	#10 counter$count = 40250;
	#10 counter$count = 40251;
	#10 counter$count = 40252;
	#10 counter$count = 40253;
	#10 counter$count = 40254;
	#10 counter$count = 40255;
	#10 counter$count = 40256;
	#10 counter$count = 40257;
	#10 counter$count = 40258;
	#10 counter$count = 40259;
	#10 counter$count = 40260;
	#10 counter$count = 40261;
	#10 counter$count = 40262;
	#10 counter$count = 40263;
	#10 counter$count = 40264;
	#10 counter$count = 40265;
	#10 counter$count = 40266;
	#10 counter$count = 40267;
	#10 counter$count = 40268;
	#10 counter$count = 40269;
	#10 counter$count = 40270;
	#10 counter$count = 40271;
	#10 counter$count = 40272;
	#10 counter$count = 40273;
	#10 counter$count = 40274;
	#10 counter$count = 40275;
	#10 counter$count = 40276;
	#10 counter$count = 40277;
	#10 counter$count = 40278;
	#10 counter$count = 40279;
	#10 counter$count = 40280;
	#10 counter$count = 40281;
	#10 counter$count = 40282;
	#10 counter$count = 40283;
	#10 counter$count = 40284;
	#10 counter$count = 40285;
	#10 counter$count = 40286;
	#10 counter$count = 40287;
	#10 counter$count = 40288;
	#10 counter$count = 40289;
	#10 counter$count = 40290;
	#10 counter$count = 40291;
	#10 counter$count = 40292;
	#10 counter$count = 40293;
	#10 counter$count = 40294;
	#10 counter$count = 40295;
	#10 counter$count = 40296;
	#10 counter$count = 40297;
	#10 counter$count = 40298;
	#10 counter$count = 40299;
	#10 counter$count = 40300;
	#10 counter$count = 40301;
	#10 counter$count = 40302;
	#10 counter$count = 40303;
	#10 counter$count = 40304;
	#10 counter$count = 40305;
	#10 counter$count = 40306;
	#10 counter$count = 40307;
	#10 counter$count = 40308;
	#10 counter$count = 40309;
	#10 counter$count = 40310;
	#10 counter$count = 40311;
	#10 counter$count = 40312;
	#10 counter$count = 40313;
	#10 counter$count = 40314;
	#10 counter$count = 40315;
	#10 counter$count = 40316;
	#10 counter$count = 40317;
	#10 counter$count = 40318;
	#10 counter$count = 40319;
	#10 counter$count = 40320;
	#10 counter$count = 40321;
	#10 counter$count = 40322;
	#10 counter$count = 40323;
	#10 counter$count = 40324;
	#10 counter$count = 40325;
	#10 counter$count = 40326;
	#10 counter$count = 40327;
	#10 counter$count = 40328;
	#10 counter$count = 40329;
	#10 counter$count = 40330;
	#10 counter$count = 40331;
	#10 counter$count = 40332;
	#10 counter$count = 40333;
	#10 counter$count = 40334;
	#10 counter$count = 40335;
	#10 counter$count = 40336;
	#10 counter$count = 40337;
	#10 counter$count = 40338;
	#10 counter$count = 40339;
	#10 counter$count = 40340;
	#10 counter$count = 40341;
	#10 counter$count = 40342;
	#10 counter$count = 40343;
	#10 counter$count = 40344;
	#10 counter$count = 40345;
	#10 counter$count = 40346;
	#10 counter$count = 40347;
	#10 counter$count = 40348;
	#10 counter$count = 40349;
	#10 counter$count = 40350;
	#10 counter$count = 40351;
	#10 counter$count = 40352;
	#10 counter$count = 40353;
	#10 counter$count = 40354;
	#10 counter$count = 40355;
	#10 counter$count = 40356;
	#10 counter$count = 40357;
	#10 counter$count = 40358;
	#10 counter$count = 40359;
	#10 counter$count = 40360;
	#10 counter$count = 40361;
	#10 counter$count = 40362;
	#10 counter$count = 40363;
	#10 counter$count = 40364;
	#10 counter$count = 40365;
	#10 counter$count = 40366;
	#10 counter$count = 40367;
	#10 counter$count = 40368;
	#10 counter$count = 40369;
	#10 counter$count = 40370;
	#10 counter$count = 40371;
	#10 counter$count = 40372;
	#10 counter$count = 40373;
	#10 counter$count = 40374;
	#10 counter$count = 40375;
	#10 counter$count = 40376;
	#10 counter$count = 40377;
	#10 counter$count = 40378;
	#10 counter$count = 40379;
	#10 counter$count = 40380;
	#10 counter$count = 40381;
	#10 counter$count = 40382;
	#10 counter$count = 40383;
	#10 counter$count = 40384;
	#10 counter$count = 40385;
	#10 counter$count = 40386;
	#10 counter$count = 40387;
	#10 counter$count = 40388;
	#10 counter$count = 40389;
	#10 counter$count = 40390;
	#10 counter$count = 40391;
	#10 counter$count = 40392;
	#10 counter$count = 40393;
	#10 counter$count = 40394;
	#10 counter$count = 40395;
	#10 counter$count = 40396;
	#10 counter$count = 40397;
	#10 counter$count = 40398;
	#10 counter$count = 40399;
	#10 counter$count = 40400;
	#10 counter$count = 40401;
	#10 counter$count = 40402;
	#10 counter$count = 40403;
	#10 counter$count = 40404;
	#10 counter$count = 40405;
	#10 counter$count = 40406;
	#10 counter$count = 40407;
	#10 counter$count = 40408;
	#10 counter$count = 40409;
	#10 counter$count = 40410;
	#10 counter$count = 40411;
	#10 counter$count = 40412;
	#10 counter$count = 40413;
	#10 counter$count = 40414;
	#10 counter$count = 40415;
	#10 counter$count = 40416;
	#10 counter$count = 40417;
	#10 counter$count = 40418;
	#10 counter$count = 40419;
	#10 counter$count = 40420;
	#10 counter$count = 40421;
	#10 counter$count = 40422;
	#10 counter$count = 40423;
	#10 counter$count = 40424;
	#10 counter$count = 40425;
	#10 counter$count = 40426;
	#10 counter$count = 40427;
	#10 counter$count = 40428;
	#10 counter$count = 40429;
	#10 counter$count = 40430;
	#10 counter$count = 40431;
	#10 counter$count = 40432;
	#10 counter$count = 40433;
	#10 counter$count = 40434;
	#10 counter$count = 40435;
	#10 counter$count = 40436;
	#10 counter$count = 40437;
	#10 counter$count = 40438;
	#10 counter$count = 40439;
	#10 counter$count = 40440;
	#10 counter$count = 40441;
	#10 counter$count = 40442;
	#10 counter$count = 40443;
	#10 counter$count = 40444;
	#10 counter$count = 40445;
	#10 counter$count = 40446;
	#10 counter$count = 40447;
	#10 counter$count = 40448;
	#10 counter$count = 40449;
	#10 counter$count = 40450;
	#10 counter$count = 40451;
	#10 counter$count = 40452;
	#10 counter$count = 40453;
	#10 counter$count = 40454;
	#10 counter$count = 40455;
	#10 counter$count = 40456;
	#10 counter$count = 40457;
	#10 counter$count = 40458;
	#10 counter$count = 40459;
	#10 counter$count = 40460;
	#10 counter$count = 40461;
	#10 counter$count = 40462;
	#10 counter$count = 40463;
	#10 counter$count = 40464;
	#10 counter$count = 40465;
	#10 counter$count = 40466;
	#10 counter$count = 40467;
	#10 counter$count = 40468;
	#10 counter$count = 40469;
	#10 counter$count = 40470;
	#10 counter$count = 40471;
	#10 counter$count = 40472;
	#10 counter$count = 40473;
	#10 counter$count = 40474;
	#10 counter$count = 40475;
	#10 counter$count = 40476;
	#10 counter$count = 40477;
	#10 counter$count = 40478;
	#10 counter$count = 40479;
	#10 counter$count = 40480;
	#10 counter$count = 40481;
	#10 counter$count = 40482;
	#10 counter$count = 40483;
	#10 counter$count = 40484;
	#10 counter$count = 40485;
	#10 counter$count = 40486;
	#10 counter$count = 40487;
	#10 counter$count = 40488;
	#10 counter$count = 40489;
	#10 counter$count = 40490;
	#10 counter$count = 40491;
	#10 counter$count = 40492;
	#10 counter$count = 40493;
	#10 counter$count = 40494;
	#10 counter$count = 40495;
	#10 counter$count = 40496;
	#10 counter$count = 40497;
	#10 counter$count = 40498;
	#10 counter$count = 40499;
	#10 counter$count = 40500;
	#10 counter$count = 40501;
	#10 counter$count = 40502;
	#10 counter$count = 40503;
	#10 counter$count = 40504;
	#10 counter$count = 40505;
	#10 counter$count = 40506;
	#10 counter$count = 40507;
	#10 counter$count = 40508;
	#10 counter$count = 40509;
	#10 counter$count = 40510;
	#10 counter$count = 40511;
	#10 counter$count = 40512;
	#10 counter$count = 40513;
	#10 counter$count = 40514;
	#10 counter$count = 40515;
	#10 counter$count = 40516;
	#10 counter$count = 40517;
	#10 counter$count = 40518;
	#10 counter$count = 40519;
	#10 counter$count = 40520;
	#10 counter$count = 40521;
	#10 counter$count = 40522;
	#10 counter$count = 40523;
	#10 counter$count = 40524;
	#10 counter$count = 40525;
	#10 counter$count = 40526;
	#10 counter$count = 40527;
	#10 counter$count = 40528;
	#10 counter$count = 40529;
	#10 counter$count = 40530;
	#10 counter$count = 40531;
	#10 counter$count = 40532;
	#10 counter$count = 40533;
	#10 counter$count = 40534;
	#10 counter$count = 40535;
	#10 counter$count = 40536;
	#10 counter$count = 40537;
	#10 counter$count = 40538;
	#10 counter$count = 40539;
	#10 counter$count = 40540;
	#10 counter$count = 40541;
	#10 counter$count = 40542;
	#10 counter$count = 40543;
	#10 counter$count = 40544;
	#10 counter$count = 40545;
	#10 counter$count = 40546;
	#10 counter$count = 40547;
	#10 counter$count = 40548;
	#10 counter$count = 40549;
	#10 counter$count = 40550;
	#10 counter$count = 40551;
	#10 counter$count = 40552;
	#10 counter$count = 40553;
	#10 counter$count = 40554;
	#10 counter$count = 40555;
	#10 counter$count = 40556;
	#10 counter$count = 40557;
	#10 counter$count = 40558;
	#10 counter$count = 40559;
	#10 counter$count = 40560;
	#10 counter$count = 40561;
	#10 counter$count = 40562;
	#10 counter$count = 40563;
	#10 counter$count = 40564;
	#10 counter$count = 40565;
	#10 counter$count = 40566;
	#10 counter$count = 40567;
	#10 counter$count = 40568;
	#10 counter$count = 40569;
	#10 counter$count = 40570;
	#10 counter$count = 40571;
	#10 counter$count = 40572;
	#10 counter$count = 40573;
	#10 counter$count = 40574;
	#10 counter$count = 40575;
	#10 counter$count = 40576;
	#10 counter$count = 40577;
	#10 counter$count = 40578;
	#10 counter$count = 40579;
	#10 counter$count = 40580;
	#10 counter$count = 40581;
	#10 counter$count = 40582;
	#10 counter$count = 40583;
	#10 counter$count = 40584;
	#10 counter$count = 40585;
	#10 counter$count = 40586;
	#10 counter$count = 40587;
	#10 counter$count = 40588;
	#10 counter$count = 40589;
	#10 counter$count = 40590;
	#10 counter$count = 40591;
	#10 counter$count = 40592;
	#10 counter$count = 40593;
	#10 counter$count = 40594;
	#10 counter$count = 40595;
	#10 counter$count = 40596;
	#10 counter$count = 40597;
	#10 counter$count = 40598;
	#10 counter$count = 40599;
	#10 counter$count = 40600;
	#10 counter$count = 40601;
	#10 counter$count = 40602;
	#10 counter$count = 40603;
	#10 counter$count = 40604;
	#10 counter$count = 40605;
	#10 counter$count = 40606;
	#10 counter$count = 40607;
	#10 counter$count = 40608;
	#10 counter$count = 40609;
	#10 counter$count = 40610;
	#10 counter$count = 40611;
	#10 counter$count = 40612;
	#10 counter$count = 40613;
	#10 counter$count = 40614;
	#10 counter$count = 40615;
	#10 counter$count = 40616;
	#10 counter$count = 40617;
	#10 counter$count = 40618;
	#10 counter$count = 40619;
	#10 counter$count = 40620;
	#10 counter$count = 40621;
	#10 counter$count = 40622;
	#10 counter$count = 40623;
	#10 counter$count = 40624;
	#10 counter$count = 40625;
	#10 counter$count = 40626;
	#10 counter$count = 40627;
	#10 counter$count = 40628;
	#10 counter$count = 40629;
	#10 counter$count = 40630;
	#10 counter$count = 40631;
	#10 counter$count = 40632;
	#10 counter$count = 40633;
	#10 counter$count = 40634;
	#10 counter$count = 40635;
	#10 counter$count = 40636;
	#10 counter$count = 40637;
	#10 counter$count = 40638;
	#10 counter$count = 40639;
	#10 counter$count = 40640;
	#10 counter$count = 40641;
	#10 counter$count = 40642;
	#10 counter$count = 40643;
	#10 counter$count = 40644;
	#10 counter$count = 40645;
	#10 counter$count = 40646;
	#10 counter$count = 40647;
	#10 counter$count = 40648;
	#10 counter$count = 40649;
	#10 counter$count = 40650;
	#10 counter$count = 40651;
	#10 counter$count = 40652;
	#10 counter$count = 40653;
	#10 counter$count = 40654;
	#10 counter$count = 40655;
	#10 counter$count = 40656;
	#10 counter$count = 40657;
	#10 counter$count = 40658;
	#10 counter$count = 40659;
	#10 counter$count = 40660;
	#10 counter$count = 40661;
	#10 counter$count = 40662;
	#10 counter$count = 40663;
	#10 counter$count = 40664;
	#10 counter$count = 40665;
	#10 counter$count = 40666;
	#10 counter$count = 40667;
	#10 counter$count = 40668;
	#10 counter$count = 40669;
	#10 counter$count = 40670;
	#10 counter$count = 40671;
	#10 counter$count = 40672;
	#10 counter$count = 40673;
	#10 counter$count = 40674;
	#10 counter$count = 40675;
	#10 counter$count = 40676;
	#10 counter$count = 40677;
	#10 counter$count = 40678;
	#10 counter$count = 40679;
	#10 counter$count = 40680;
	#10 counter$count = 40681;
	#10 counter$count = 40682;
	#10 counter$count = 40683;
	#10 counter$count = 40684;
	#10 counter$count = 40685;
	#10 counter$count = 40686;
	#10 counter$count = 40687;
	#10 counter$count = 40688;
	#10 counter$count = 40689;
	#10 counter$count = 40690;
	#10 counter$count = 40691;
	#10 counter$count = 40692;
	#10 counter$count = 40693;
	#10 counter$count = 40694;
	#10 counter$count = 40695;
	#10 counter$count = 40696;
	#10 counter$count = 40697;
	#10 counter$count = 40698;
	#10 counter$count = 40699;
	#10 counter$count = 40700;
	#10 counter$count = 40701;
	#10 counter$count = 40702;
	#10 counter$count = 40703;
	#10 counter$count = 40704;
	#10 counter$count = 40705;
	#10 counter$count = 40706;
	#10 counter$count = 40707;
	#10 counter$count = 40708;
	#10 counter$count = 40709;
	#10 counter$count = 40710;
	#10 counter$count = 40711;
	#10 counter$count = 40712;
	#10 counter$count = 40713;
	#10 counter$count = 40714;
	#10 counter$count = 40715;
	#10 counter$count = 40716;
	#10 counter$count = 40717;
	#10 counter$count = 40718;
	#10 counter$count = 40719;
	#10 counter$count = 40720;
	#10 counter$count = 40721;
	#10 counter$count = 40722;
	#10 counter$count = 40723;
	#10 counter$count = 40724;
	#10 counter$count = 40725;
	#10 counter$count = 40726;
	#10 counter$count = 40727;
	#10 counter$count = 40728;
	#10 counter$count = 40729;
	#10 counter$count = 40730;
	#10 counter$count = 40731;
	#10 counter$count = 40732;
	#10 counter$count = 40733;
	#10 counter$count = 40734;
	#10 counter$count = 40735;
	#10 counter$count = 40736;
	#10 counter$count = 40737;
	#10 counter$count = 40738;
	#10 counter$count = 40739;
	#10 counter$count = 40740;
	#10 counter$count = 40741;
	#10 counter$count = 40742;
	#10 counter$count = 40743;
	#10 counter$count = 40744;
	#10 counter$count = 40745;
	#10 counter$count = 40746;
	#10 counter$count = 40747;
	#10 counter$count = 40748;
	#10 counter$count = 40749;
	#10 counter$count = 40750;
	#10 counter$count = 40751;
	#10 counter$count = 40752;
	#10 counter$count = 40753;
	#10 counter$count = 40754;
	#10 counter$count = 40755;
	#10 counter$count = 40756;
	#10 counter$count = 40757;
	#10 counter$count = 40758;
	#10 counter$count = 40759;
	#10 counter$count = 40760;
	#10 counter$count = 40761;
	#10 counter$count = 40762;
	#10 counter$count = 40763;
	#10 counter$count = 40764;
	#10 counter$count = 40765;
	#10 counter$count = 40766;
	#10 counter$count = 40767;
	#10 counter$count = 40768;
	#10 counter$count = 40769;
	#10 counter$count = 40770;
	#10 counter$count = 40771;
	#10 counter$count = 40772;
	#10 counter$count = 40773;
	#10 counter$count = 40774;
	#10 counter$count = 40775;
	#10 counter$count = 40776;
	#10 counter$count = 40777;
	#10 counter$count = 40778;
	#10 counter$count = 40779;
	#10 counter$count = 40780;
	#10 counter$count = 40781;
	#10 counter$count = 40782;
	#10 counter$count = 40783;
	#10 counter$count = 40784;
	#10 counter$count = 40785;
	#10 counter$count = 40786;
	#10 counter$count = 40787;
	#10 counter$count = 40788;
	#10 counter$count = 40789;
	#10 counter$count = 40790;
	#10 counter$count = 40791;
	#10 counter$count = 40792;
	#10 counter$count = 40793;
	#10 counter$count = 40794;
	#10 counter$count = 40795;
	#10 counter$count = 40796;
	#10 counter$count = 40797;
	#10 counter$count = 40798;
	#10 counter$count = 40799;
	#10 counter$count = 40800;
	#10 counter$count = 40801;
	#10 counter$count = 40802;
	#10 counter$count = 40803;
	#10 counter$count = 40804;
	#10 counter$count = 40805;
	#10 counter$count = 40806;
	#10 counter$count = 40807;
	#10 counter$count = 40808;
	#10 counter$count = 40809;
	#10 counter$count = 40810;
	#10 counter$count = 40811;
	#10 counter$count = 40812;
	#10 counter$count = 40813;
	#10 counter$count = 40814;
	#10 counter$count = 40815;
	#10 counter$count = 40816;
	#10 counter$count = 40817;
	#10 counter$count = 40818;
	#10 counter$count = 40819;
	#10 counter$count = 40820;
	#10 counter$count = 40821;
	#10 counter$count = 40822;
	#10 counter$count = 40823;
	#10 counter$count = 40824;
	#10 counter$count = 40825;
	#10 counter$count = 40826;
	#10 counter$count = 40827;
	#10 counter$count = 40828;
	#10 counter$count = 40829;
	#10 counter$count = 40830;
	#10 counter$count = 40831;
	#10 counter$count = 40832;
	#10 counter$count = 40833;
	#10 counter$count = 40834;
	#10 counter$count = 40835;
	#10 counter$count = 40836;
	#10 counter$count = 40837;
	#10 counter$count = 40838;
	#10 counter$count = 40839;
	#10 counter$count = 40840;
	#10 counter$count = 40841;
	#10 counter$count = 40842;
	#10 counter$count = 40843;
	#10 counter$count = 40844;
	#10 counter$count = 40845;
	#10 counter$count = 40846;
	#10 counter$count = 40847;
	#10 counter$count = 40848;
	#10 counter$count = 40849;
	#10 counter$count = 40850;
	#10 counter$count = 40851;
	#10 counter$count = 40852;
	#10 counter$count = 40853;
	#10 counter$count = 40854;
	#10 counter$count = 40855;
	#10 counter$count = 40856;
	#10 counter$count = 40857;
	#10 counter$count = 40858;
	#10 counter$count = 40859;
	#10 counter$count = 40860;
	#10 counter$count = 40861;
	#10 counter$count = 40862;
	#10 counter$count = 40863;
	#10 counter$count = 40864;
	#10 counter$count = 40865;
	#10 counter$count = 40866;
	#10 counter$count = 40867;
	#10 counter$count = 40868;
	#10 counter$count = 40869;
	#10 counter$count = 40870;
	#10 counter$count = 40871;
	#10 counter$count = 40872;
	#10 counter$count = 40873;
	#10 counter$count = 40874;
	#10 counter$count = 40875;
	#10 counter$count = 40876;
	#10 counter$count = 40877;
	#10 counter$count = 40878;
	#10 counter$count = 40879;
	#10 counter$count = 40880;
	#10 counter$count = 40881;
	#10 counter$count = 40882;
	#10 counter$count = 40883;
	#10 counter$count = 40884;
	#10 counter$count = 40885;
	#10 counter$count = 40886;
	#10 counter$count = 40887;
	#10 counter$count = 40888;
	#10 counter$count = 40889;
	#10 counter$count = 40890;
	#10 counter$count = 40891;
	#10 counter$count = 40892;
	#10 counter$count = 40893;
	#10 counter$count = 40894;
	#10 counter$count = 40895;
	#10 counter$count = 40896;
	#10 counter$count = 40897;
	#10 counter$count = 40898;
	#10 counter$count = 40899;
	#10 counter$count = 40900;
	#10 counter$count = 40901;
	#10 counter$count = 40902;
	#10 counter$count = 40903;
	#10 counter$count = 40904;
	#10 counter$count = 40905;
	#10 counter$count = 40906;
	#10 counter$count = 40907;
	#10 counter$count = 40908;
	#10 counter$count = 40909;
	#10 counter$count = 40910;
	#10 counter$count = 40911;
	#10 counter$count = 40912;
	#10 counter$count = 40913;
	#10 counter$count = 40914;
	#10 counter$count = 40915;
	#10 counter$count = 40916;
	#10 counter$count = 40917;
	#10 counter$count = 40918;
	#10 counter$count = 40919;
	#10 counter$count = 40920;
	#10 counter$count = 40921;
	#10 counter$count = 40922;
	#10 counter$count = 40923;
	#10 counter$count = 40924;
	#10 counter$count = 40925;
	#10 counter$count = 40926;
	#10 counter$count = 40927;
	#10 counter$count = 40928;
	#10 counter$count = 40929;
	#10 counter$count = 40930;
	#10 counter$count = 40931;
	#10 counter$count = 40932;
	#10 counter$count = 40933;
	#10 counter$count = 40934;
	#10 counter$count = 40935;
	#10 counter$count = 40936;
	#10 counter$count = 40937;
	#10 counter$count = 40938;
	#10 counter$count = 40939;
	#10 counter$count = 40940;
	#10 counter$count = 40941;
	#10 counter$count = 40942;
	#10 counter$count = 40943;
	#10 counter$count = 40944;
	#10 counter$count = 40945;
	#10 counter$count = 40946;
	#10 counter$count = 40947;
	#10 counter$count = 40948;
	#10 counter$count = 40949;
	#10 counter$count = 40950;
	#10 counter$count = 40951;
	#10 counter$count = 40952;
	#10 counter$count = 40953;
	#10 counter$count = 40954;
	#10 counter$count = 40955;
	#10 counter$count = 40956;
	#10 counter$count = 40957;
	#10 counter$count = 40958;
	#10 counter$count = 40959;
	#10 counter$count = 40960;
	#10 counter$count = 40961;
	#10 counter$count = 40962;
	#10 counter$count = 40963;
	#10 counter$count = 40964;
	#10 counter$count = 40965;
	#10 counter$count = 40966;
	#10 counter$count = 40967;
	#10 counter$count = 40968;
	#10 counter$count = 40969;
	#10 counter$count = 40970;
	#10 counter$count = 40971;
	#10 counter$count = 40972;
	#10 counter$count = 40973;
	#10 counter$count = 40974;
	#10 counter$count = 40975;
	#10 counter$count = 40976;
	#10 counter$count = 40977;
	#10 counter$count = 40978;
	#10 counter$count = 40979;
	#10 counter$count = 40980;
	#10 counter$count = 40981;
	#10 counter$count = 40982;
	#10 counter$count = 40983;
	#10 counter$count = 40984;
	#10 counter$count = 40985;
	#10 counter$count = 40986;
	#10 counter$count = 40987;
	#10 counter$count = 40988;
	#10 counter$count = 40989;
	#10 counter$count = 40990;
	#10 counter$count = 40991;
	#10 counter$count = 40992;
	#10 counter$count = 40993;
	#10 counter$count = 40994;
	#10 counter$count = 40995;
	#10 counter$count = 40996;
	#10 counter$count = 40997;
	#10 counter$count = 40998;
	#10 counter$count = 40999;
	#10 counter$count = 41000;
	#10 counter$count = 41001;
	#10 counter$count = 41002;
	#10 counter$count = 41003;
	#10 counter$count = 41004;
	#10 counter$count = 41005;
	#10 counter$count = 41006;
	#10 counter$count = 41007;
	#10 counter$count = 41008;
	#10 counter$count = 41009;
	#10 counter$count = 41010;
	#10 counter$count = 41011;
	#10 counter$count = 41012;
	#10 counter$count = 41013;
	#10 counter$count = 41014;
	#10 counter$count = 41015;
	#10 counter$count = 41016;
	#10 counter$count = 41017;
	#10 counter$count = 41018;
	#10 counter$count = 41019;
	#10 counter$count = 41020;
	#10 counter$count = 41021;
	#10 counter$count = 41022;
	#10 counter$count = 41023;
	#10 counter$count = 41024;
	#10 counter$count = 41025;
	#10 counter$count = 41026;
	#10 counter$count = 41027;
	#10 counter$count = 41028;
	#10 counter$count = 41029;
	#10 counter$count = 41030;
	#10 counter$count = 41031;
	#10 counter$count = 41032;
	#10 counter$count = 41033;
	#10 counter$count = 41034;
	#10 counter$count = 41035;
	#10 counter$count = 41036;
	#10 counter$count = 41037;
	#10 counter$count = 41038;
	#10 counter$count = 41039;
	#10 counter$count = 41040;
	#10 counter$count = 41041;
	#10 counter$count = 41042;
	#10 counter$count = 41043;
	#10 counter$count = 41044;
	#10 counter$count = 41045;
	#10 counter$count = 41046;
	#10 counter$count = 41047;
	#10 counter$count = 41048;
	#10 counter$count = 41049;
	#10 counter$count = 41050;
	#10 counter$count = 41051;
	#10 counter$count = 41052;
	#10 counter$count = 41053;
	#10 counter$count = 41054;
	#10 counter$count = 41055;
	#10 counter$count = 41056;
	#10 counter$count = 41057;
	#10 counter$count = 41058;
	#10 counter$count = 41059;
	#10 counter$count = 41060;
	#10 counter$count = 41061;
	#10 counter$count = 41062;
	#10 counter$count = 41063;
	#10 counter$count = 41064;
	#10 counter$count = 41065;
	#10 counter$count = 41066;
	#10 counter$count = 41067;
	#10 counter$count = 41068;
	#10 counter$count = 41069;
	#10 counter$count = 41070;
	#10 counter$count = 41071;
	#10 counter$count = 41072;
	#10 counter$count = 41073;
	#10 counter$count = 41074;
	#10 counter$count = 41075;
	#10 counter$count = 41076;
	#10 counter$count = 41077;
	#10 counter$count = 41078;
	#10 counter$count = 41079;
	#10 counter$count = 41080;
	#10 counter$count = 41081;
	#10 counter$count = 41082;
	#10 counter$count = 41083;
	#10 counter$count = 41084;
	#10 counter$count = 41085;
	#10 counter$count = 41086;
	#10 counter$count = 41087;
	#10 counter$count = 41088;
	#10 counter$count = 41089;
	#10 counter$count = 41090;
	#10 counter$count = 41091;
	#10 counter$count = 41092;
	#10 counter$count = 41093;
	#10 counter$count = 41094;
	#10 counter$count = 41095;
	#10 counter$count = 41096;
	#10 counter$count = 41097;
	#10 counter$count = 41098;
	#10 counter$count = 41099;
	#10 counter$count = 41100;
	#10 counter$count = 41101;
	#10 counter$count = 41102;
	#10 counter$count = 41103;
	#10 counter$count = 41104;
	#10 counter$count = 41105;
	#10 counter$count = 41106;
	#10 counter$count = 41107;
	#10 counter$count = 41108;
	#10 counter$count = 41109;
	#10 counter$count = 41110;
	#10 counter$count = 41111;
	#10 counter$count = 41112;
	#10 counter$count = 41113;
	#10 counter$count = 41114;
	#10 counter$count = 41115;
	#10 counter$count = 41116;
	#10 counter$count = 41117;
	#10 counter$count = 41118;
	#10 counter$count = 41119;
	#10 counter$count = 41120;
	#10 counter$count = 41121;
	#10 counter$count = 41122;
	#10 counter$count = 41123;
	#10 counter$count = 41124;
	#10 counter$count = 41125;
	#10 counter$count = 41126;
	#10 counter$count = 41127;
	#10 counter$count = 41128;
	#10 counter$count = 41129;
	#10 counter$count = 41130;
	#10 counter$count = 41131;
	#10 counter$count = 41132;
	#10 counter$count = 41133;
	#10 counter$count = 41134;
	#10 counter$count = 41135;
	#10 counter$count = 41136;
	#10 counter$count = 41137;
	#10 counter$count = 41138;
	#10 counter$count = 41139;
	#10 counter$count = 41140;
	#10 counter$count = 41141;
	#10 counter$count = 41142;
	#10 counter$count = 41143;
	#10 counter$count = 41144;
	#10 counter$count = 41145;
	#10 counter$count = 41146;
	#10 counter$count = 41147;
	#10 counter$count = 41148;
	#10 counter$count = 41149;
	#10 counter$count = 41150;
	#10 counter$count = 41151;
	#10 counter$count = 41152;
	#10 counter$count = 41153;
	#10 counter$count = 41154;
	#10 counter$count = 41155;
	#10 counter$count = 41156;
	#10 counter$count = 41157;
	#10 counter$count = 41158;
	#10 counter$count = 41159;
	#10 counter$count = 41160;
	#10 counter$count = 41161;
	#10 counter$count = 41162;
	#10 counter$count = 41163;
	#10 counter$count = 41164;
	#10 counter$count = 41165;
	#10 counter$count = 41166;
	#10 counter$count = 41167;
	#10 counter$count = 41168;
	#10 counter$count = 41169;
	#10 counter$count = 41170;
	#10 counter$count = 41171;
	#10 counter$count = 41172;
	#10 counter$count = 41173;
	#10 counter$count = 41174;
	#10 counter$count = 41175;
	#10 counter$count = 41176;
	#10 counter$count = 41177;
	#10 counter$count = 41178;
	#10 counter$count = 41179;
	#10 counter$count = 41180;
	#10 counter$count = 41181;
	#10 counter$count = 41182;
	#10 counter$count = 41183;
	#10 counter$count = 41184;
	#10 counter$count = 41185;
	#10 counter$count = 41186;
	#10 counter$count = 41187;
	#10 counter$count = 41188;
	#10 counter$count = 41189;
	#10 counter$count = 41190;
	#10 counter$count = 41191;
	#10 counter$count = 41192;
	#10 counter$count = 41193;
	#10 counter$count = 41194;
	#10 counter$count = 41195;
	#10 counter$count = 41196;
	#10 counter$count = 41197;
	#10 counter$count = 41198;
	#10 counter$count = 41199;
	#10 counter$count = 41200;
	#10 counter$count = 41201;
	#10 counter$count = 41202;
	#10 counter$count = 41203;
	#10 counter$count = 41204;
	#10 counter$count = 41205;
	#10 counter$count = 41206;
	#10 counter$count = 41207;
	#10 counter$count = 41208;
	#10 counter$count = 41209;
	#10 counter$count = 41210;
	#10 counter$count = 41211;
	#10 counter$count = 41212;
	#10 counter$count = 41213;
	#10 counter$count = 41214;
	#10 counter$count = 41215;
	#10 counter$count = 41216;
	#10 counter$count = 41217;
	#10 counter$count = 41218;
	#10 counter$count = 41219;
	#10 counter$count = 41220;
	#10 counter$count = 41221;
	#10 counter$count = 41222;
	#10 counter$count = 41223;
	#10 counter$count = 41224;
	#10 counter$count = 41225;
	#10 counter$count = 41226;
	#10 counter$count = 41227;
	#10 counter$count = 41228;
	#10 counter$count = 41229;
	#10 counter$count = 41230;
	#10 counter$count = 41231;
	#10 counter$count = 41232;
	#10 counter$count = 41233;
	#10 counter$count = 41234;
	#10 counter$count = 41235;
	#10 counter$count = 41236;
	#10 counter$count = 41237;
	#10 counter$count = 41238;
	#10 counter$count = 41239;
	#10 counter$count = 41240;
	#10 counter$count = 41241;
	#10 counter$count = 41242;
	#10 counter$count = 41243;
	#10 counter$count = 41244;
	#10 counter$count = 41245;
	#10 counter$count = 41246;
	#10 counter$count = 41247;
	#10 counter$count = 41248;
	#10 counter$count = 41249;
	#10 counter$count = 41250;
	#10 counter$count = 41251;
	#10 counter$count = 41252;
	#10 counter$count = 41253;
	#10 counter$count = 41254;
	#10 counter$count = 41255;
	#10 counter$count = 41256;
	#10 counter$count = 41257;
	#10 counter$count = 41258;
	#10 counter$count = 41259;
	#10 counter$count = 41260;
	#10 counter$count = 41261;
	#10 counter$count = 41262;
	#10 counter$count = 41263;
	#10 counter$count = 41264;
	#10 counter$count = 41265;
	#10 counter$count = 41266;
	#10 counter$count = 41267;
	#10 counter$count = 41268;
	#10 counter$count = 41269;
	#10 counter$count = 41270;
	#10 counter$count = 41271;
	#10 counter$count = 41272;
	#10 counter$count = 41273;
	#10 counter$count = 41274;
	#10 counter$count = 41275;
	#10 counter$count = 41276;
	#10 counter$count = 41277;
	#10 counter$count = 41278;
	#10 counter$count = 41279;
	#10 counter$count = 41280;
	#10 counter$count = 41281;
	#10 counter$count = 41282;
	#10 counter$count = 41283;
	#10 counter$count = 41284;
	#10 counter$count = 41285;
	#10 counter$count = 41286;
	#10 counter$count = 41287;
	#10 counter$count = 41288;
	#10 counter$count = 41289;
	#10 counter$count = 41290;
	#10 counter$count = 41291;
	#10 counter$count = 41292;
	#10 counter$count = 41293;
	#10 counter$count = 41294;
	#10 counter$count = 41295;
	#10 counter$count = 41296;
	#10 counter$count = 41297;
	#10 counter$count = 41298;
	#10 counter$count = 41299;
	#10 counter$count = 41300;
	#10 counter$count = 41301;
	#10 counter$count = 41302;
	#10 counter$count = 41303;
	#10 counter$count = 41304;
	#10 counter$count = 41305;
	#10 counter$count = 41306;
	#10 counter$count = 41307;
	#10 counter$count = 41308;
	#10 counter$count = 41309;
	#10 counter$count = 41310;
	#10 counter$count = 41311;
	#10 counter$count = 41312;
	#10 counter$count = 41313;
	#10 counter$count = 41314;
	#10 counter$count = 41315;
	#10 counter$count = 41316;
	#10 counter$count = 41317;
	#10 counter$count = 41318;
	#10 counter$count = 41319;
	#10 counter$count = 41320;
	#10 counter$count = 41321;
	#10 counter$count = 41322;
	#10 counter$count = 41323;
	#10 counter$count = 41324;
	#10 counter$count = 41325;
	#10 counter$count = 41326;
	#10 counter$count = 41327;
	#10 counter$count = 41328;
	#10 counter$count = 41329;
	#10 counter$count = 41330;
	#10 counter$count = 41331;
	#10 counter$count = 41332;
	#10 counter$count = 41333;
	#10 counter$count = 41334;
	#10 counter$count = 41335;
	#10 counter$count = 41336;
	#10 counter$count = 41337;
	#10 counter$count = 41338;
	#10 counter$count = 41339;
	#10 counter$count = 41340;
	#10 counter$count = 41341;
	#10 counter$count = 41342;
	#10 counter$count = 41343;
	#10 counter$count = 41344;
	#10 counter$count = 41345;
	#10 counter$count = 41346;
	#10 counter$count = 41347;
	#10 counter$count = 41348;
	#10 counter$count = 41349;
	#10 counter$count = 41350;
	#10 counter$count = 41351;
	#10 counter$count = 41352;
	#10 counter$count = 41353;
	#10 counter$count = 41354;
	#10 counter$count = 41355;
	#10 counter$count = 41356;
	#10 counter$count = 41357;
	#10 counter$count = 41358;
	#10 counter$count = 41359;
	#10 counter$count = 41360;
	#10 counter$count = 41361;
	#10 counter$count = 41362;
	#10 counter$count = 41363;
	#10 counter$count = 41364;
	#10 counter$count = 41365;
	#10 counter$count = 41366;
	#10 counter$count = 41367;
	#10 counter$count = 41368;
	#10 counter$count = 41369;
	#10 counter$count = 41370;
	#10 counter$count = 41371;
	#10 counter$count = 41372;
	#10 counter$count = 41373;
	#10 counter$count = 41374;
	#10 counter$count = 41375;
	#10 counter$count = 41376;
	#10 counter$count = 41377;
	#10 counter$count = 41378;
	#10 counter$count = 41379;
	#10 counter$count = 41380;
	#10 counter$count = 41381;
	#10 counter$count = 41382;
	#10 counter$count = 41383;
	#10 counter$count = 41384;
	#10 counter$count = 41385;
	#10 counter$count = 41386;
	#10 counter$count = 41387;
	#10 counter$count = 41388;
	#10 counter$count = 41389;
	#10 counter$count = 41390;
	#10 counter$count = 41391;
	#10 counter$count = 41392;
	#10 counter$count = 41393;
	#10 counter$count = 41394;
	#10 counter$count = 41395;
	#10 counter$count = 41396;
	#10 counter$count = 41397;
	#10 counter$count = 41398;
	#10 counter$count = 41399;
	#10 counter$count = 41400;
	#10 counter$count = 41401;
	#10 counter$count = 41402;
	#10 counter$count = 41403;
	#10 counter$count = 41404;
	#10 counter$count = 41405;
	#10 counter$count = 41406;
	#10 counter$count = 41407;
	#10 counter$count = 41408;
	#10 counter$count = 41409;
	#10 counter$count = 41410;
	#10 counter$count = 41411;
	#10 counter$count = 41412;
	#10 counter$count = 41413;
	#10 counter$count = 41414;
	#10 counter$count = 41415;
	#10 counter$count = 41416;
	#10 counter$count = 41417;
	#10 counter$count = 41418;
	#10 counter$count = 41419;
	#10 counter$count = 41420;
	#10 counter$count = 41421;
	#10 counter$count = 41422;
	#10 counter$count = 41423;
	#10 counter$count = 41424;
	#10 counter$count = 41425;
	#10 counter$count = 41426;
	#10 counter$count = 41427;
	#10 counter$count = 41428;
	#10 counter$count = 41429;
	#10 counter$count = 41430;
	#10 counter$count = 41431;
	#10 counter$count = 41432;
	#10 counter$count = 41433;
	#10 counter$count = 41434;
	#10 counter$count = 41435;
	#10 counter$count = 41436;
	#10 counter$count = 41437;
	#10 counter$count = 41438;
	#10 counter$count = 41439;
	#10 counter$count = 41440;
	#10 counter$count = 41441;
	#10 counter$count = 41442;
	#10 counter$count = 41443;
	#10 counter$count = 41444;
	#10 counter$count = 41445;
	#10 counter$count = 41446;
	#10 counter$count = 41447;
	#10 counter$count = 41448;
	#10 counter$count = 41449;
	#10 counter$count = 41450;
	#10 counter$count = 41451;
	#10 counter$count = 41452;
	#10 counter$count = 41453;
	#10 counter$count = 41454;
	#10 counter$count = 41455;
	#10 counter$count = 41456;
	#10 counter$count = 41457;
	#10 counter$count = 41458;
	#10 counter$count = 41459;
	#10 counter$count = 41460;
	#10 counter$count = 41461;
	#10 counter$count = 41462;
	#10 counter$count = 41463;
	#10 counter$count = 41464;
	#10 counter$count = 41465;
	#10 counter$count = 41466;
	#10 counter$count = 41467;
	#10 counter$count = 41468;
	#10 counter$count = 41469;
	#10 counter$count = 41470;
	#10 counter$count = 41471;
	#10 counter$count = 41472;
	#10 counter$count = 41473;
	#10 counter$count = 41474;
	#10 counter$count = 41475;
	#10 counter$count = 41476;
	#10 counter$count = 41477;
	#10 counter$count = 41478;
	#10 counter$count = 41479;
	#10 counter$count = 41480;
	#10 counter$count = 41481;
	#10 counter$count = 41482;
	#10 counter$count = 41483;
	#10 counter$count = 41484;
	#10 counter$count = 41485;
	#10 counter$count = 41486;
	#10 counter$count = 41487;
	#10 counter$count = 41488;
	#10 counter$count = 41489;
	#10 counter$count = 41490;
	#10 counter$count = 41491;
	#10 counter$count = 41492;
	#10 counter$count = 41493;
	#10 counter$count = 41494;
	#10 counter$count = 41495;
	#10 counter$count = 41496;
	#10 counter$count = 41497;
	#10 counter$count = 41498;
	#10 counter$count = 41499;
	#10 counter$count = 41500;
	#10 counter$count = 41501;
	#10 counter$count = 41502;
	#10 counter$count = 41503;
	#10 counter$count = 41504;
	#10 counter$count = 41505;
	#10 counter$count = 41506;
	#10 counter$count = 41507;
	#10 counter$count = 41508;
	#10 counter$count = 41509;
	#10 counter$count = 41510;
	#10 counter$count = 41511;
	#10 counter$count = 41512;
	#10 counter$count = 41513;
	#10 counter$count = 41514;
	#10 counter$count = 41515;
	#10 counter$count = 41516;
	#10 counter$count = 41517;
	#10 counter$count = 41518;
	#10 counter$count = 41519;
	#10 counter$count = 41520;
	#10 counter$count = 41521;
	#10 counter$count = 41522;
	#10 counter$count = 41523;
	#10 counter$count = 41524;
	#10 counter$count = 41525;
	#10 counter$count = 41526;
	#10 counter$count = 41527;
	#10 counter$count = 41528;
	#10 counter$count = 41529;
	#10 counter$count = 41530;
	#10 counter$count = 41531;
	#10 counter$count = 41532;
	#10 counter$count = 41533;
	#10 counter$count = 41534;
	#10 counter$count = 41535;
	#10 counter$count = 41536;
	#10 counter$count = 41537;
	#10 counter$count = 41538;
	#10 counter$count = 41539;
	#10 counter$count = 41540;
	#10 counter$count = 41541;
	#10 counter$count = 41542;
	#10 counter$count = 41543;
	#10 counter$count = 41544;
	#10 counter$count = 41545;
	#10 counter$count = 41546;
	#10 counter$count = 41547;
	#10 counter$count = 41548;
	#10 counter$count = 41549;
	#10 counter$count = 41550;
	#10 counter$count = 41551;
	#10 counter$count = 41552;
	#10 counter$count = 41553;
	#10 counter$count = 41554;
	#10 counter$count = 41555;
	#10 counter$count = 41556;
	#10 counter$count = 41557;
	#10 counter$count = 41558;
	#10 counter$count = 41559;
	#10 counter$count = 41560;
	#10 counter$count = 41561;
	#10 counter$count = 41562;
	#10 counter$count = 41563;
	#10 counter$count = 41564;
	#10 counter$count = 41565;
	#10 counter$count = 41566;
	#10 counter$count = 41567;
	#10 counter$count = 41568;
	#10 counter$count = 41569;
	#10 counter$count = 41570;
	#10 counter$count = 41571;
	#10 counter$count = 41572;
	#10 counter$count = 41573;
	#10 counter$count = 41574;
	#10 counter$count = 41575;
	#10 counter$count = 41576;
	#10 counter$count = 41577;
	#10 counter$count = 41578;
	#10 counter$count = 41579;
	#10 counter$count = 41580;
	#10 counter$count = 41581;
	#10 counter$count = 41582;
	#10 counter$count = 41583;
	#10 counter$count = 41584;
	#10 counter$count = 41585;
	#10 counter$count = 41586;
	#10 counter$count = 41587;
	#10 counter$count = 41588;
	#10 counter$count = 41589;
	#10 counter$count = 41590;
	#10 counter$count = 41591;
	#10 counter$count = 41592;
	#10 counter$count = 41593;
	#10 counter$count = 41594;
	#10 counter$count = 41595;
	#10 counter$count = 41596;
	#10 counter$count = 41597;
	#10 counter$count = 41598;
	#10 counter$count = 41599;
	#10 counter$count = 41600;
	#10 counter$count = 41601;
	#10 counter$count = 41602;
	#10 counter$count = 41603;
	#10 counter$count = 41604;
	#10 counter$count = 41605;
	#10 counter$count = 41606;
	#10 counter$count = 41607;
	#10 counter$count = 41608;
	#10 counter$count = 41609;
	#10 counter$count = 41610;
	#10 counter$count = 41611;
	#10 counter$count = 41612;
	#10 counter$count = 41613;
	#10 counter$count = 41614;
	#10 counter$count = 41615;
	#10 counter$count = 41616;
	#10 counter$count = 41617;
	#10 counter$count = 41618;
	#10 counter$count = 41619;
	#10 counter$count = 41620;
	#10 counter$count = 41621;
	#10 counter$count = 41622;
	#10 counter$count = 41623;
	#10 counter$count = 41624;
	#10 counter$count = 41625;
	#10 counter$count = 41626;
	#10 counter$count = 41627;
	#10 counter$count = 41628;
	#10 counter$count = 41629;
	#10 counter$count = 41630;
	#10 counter$count = 41631;
	#10 counter$count = 41632;
	#10 counter$count = 41633;
	#10 counter$count = 41634;
	#10 counter$count = 41635;
	#10 counter$count = 41636;
	#10 counter$count = 41637;
	#10 counter$count = 41638;
	#10 counter$count = 41639;
	#10 counter$count = 41640;
	#10 counter$count = 41641;
	#10 counter$count = 41642;
	#10 counter$count = 41643;
	#10 counter$count = 41644;
	#10 counter$count = 41645;
	#10 counter$count = 41646;
	#10 counter$count = 41647;
	#10 counter$count = 41648;
	#10 counter$count = 41649;
	#10 counter$count = 41650;
	#10 counter$count = 41651;
	#10 counter$count = 41652;
	#10 counter$count = 41653;
	#10 counter$count = 41654;
	#10 counter$count = 41655;
	#10 counter$count = 41656;
	#10 counter$count = 41657;
	#10 counter$count = 41658;
	#10 counter$count = 41659;
	#10 counter$count = 41660;
	#10 counter$count = 41661;
	#10 counter$count = 41662;
	#10 counter$count = 41663;
	#10 counter$count = 41664;
	#10 counter$count = 41665;
	#10 counter$count = 41666;
	#10 counter$count = 41667;
	#10 counter$count = 41668;
	#10 counter$count = 41669;
	#10 counter$count = 41670;
	#10 counter$count = 41671;
	#10 counter$count = 41672;
	#10 counter$count = 41673;
	#10 counter$count = 41674;
	#10 counter$count = 41675;
	#10 counter$count = 41676;
	#10 counter$count = 41677;
	#10 counter$count = 41678;
	#10 counter$count = 41679;
	#10 counter$count = 41680;
	#10 counter$count = 41681;
	#10 counter$count = 41682;
	#10 counter$count = 41683;
	#10 counter$count = 41684;
	#10 counter$count = 41685;
	#10 counter$count = 41686;
	#10 counter$count = 41687;
	#10 counter$count = 41688;
	#10 counter$count = 41689;
	#10 counter$count = 41690;
	#10 counter$count = 41691;
	#10 counter$count = 41692;
	#10 counter$count = 41693;
	#10 counter$count = 41694;
	#10 counter$count = 41695;
	#10 counter$count = 41696;
	#10 counter$count = 41697;
	#10 counter$count = 41698;
	#10 counter$count = 41699;
	#10 counter$count = 41700;
	#10 counter$count = 41701;
	#10 counter$count = 41702;
	#10 counter$count = 41703;
	#10 counter$count = 41704;
	#10 counter$count = 41705;
	#10 counter$count = 41706;
	#10 counter$count = 41707;
	#10 counter$count = 41708;
	#10 counter$count = 41709;
	#10 counter$count = 41710;
	#10 counter$count = 41711;
	#10 counter$count = 41712;
	#10 counter$count = 41713;
	#10 counter$count = 41714;
	#10 counter$count = 41715;
	#10 counter$count = 41716;
	#10 counter$count = 41717;
	#10 counter$count = 41718;
	#10 counter$count = 41719;
	#10 counter$count = 41720;
	#10 counter$count = 41721;
	#10 counter$count = 41722;
	#10 counter$count = 41723;
	#10 counter$count = 41724;
	#10 counter$count = 41725;
	#10 counter$count = 41726;
	#10 counter$count = 41727;
	#10 counter$count = 41728;
	#10 counter$count = 41729;
	#10 counter$count = 41730;
	#10 counter$count = 41731;
	#10 counter$count = 41732;
	#10 counter$count = 41733;
	#10 counter$count = 41734;
	#10 counter$count = 41735;
	#10 counter$count = 41736;
	#10 counter$count = 41737;
	#10 counter$count = 41738;
	#10 counter$count = 41739;
	#10 counter$count = 41740;
	#10 counter$count = 41741;
	#10 counter$count = 41742;
	#10 counter$count = 41743;
	#10 counter$count = 41744;
	#10 counter$count = 41745;
	#10 counter$count = 41746;
	#10 counter$count = 41747;
	#10 counter$count = 41748;
	#10 counter$count = 41749;
	#10 counter$count = 41750;
	#10 counter$count = 41751;
	#10 counter$count = 41752;
	#10 counter$count = 41753;
	#10 counter$count = 41754;
	#10 counter$count = 41755;
	#10 counter$count = 41756;
	#10 counter$count = 41757;
	#10 counter$count = 41758;
	#10 counter$count = 41759;
	#10 counter$count = 41760;
	#10 counter$count = 41761;
	#10 counter$count = 41762;
	#10 counter$count = 41763;
	#10 counter$count = 41764;
	#10 counter$count = 41765;
	#10 counter$count = 41766;
	#10 counter$count = 41767;
	#10 counter$count = 41768;
	#10 counter$count = 41769;
	#10 counter$count = 41770;
	#10 counter$count = 41771;
	#10 counter$count = 41772;
	#10 counter$count = 41773;
	#10 counter$count = 41774;
	#10 counter$count = 41775;
	#10 counter$count = 41776;
	#10 counter$count = 41777;
	#10 counter$count = 41778;
	#10 counter$count = 41779;
	#10 counter$count = 41780;
	#10 counter$count = 41781;
	#10 counter$count = 41782;
	#10 counter$count = 41783;
	#10 counter$count = 41784;
	#10 counter$count = 41785;
	#10 counter$count = 41786;
	#10 counter$count = 41787;
	#10 counter$count = 41788;
	#10 counter$count = 41789;
	#10 counter$count = 41790;
	#10 counter$count = 41791;
	#10 counter$count = 41792;
	#10 counter$count = 41793;
	#10 counter$count = 41794;
	#10 counter$count = 41795;
	#10 counter$count = 41796;
	#10 counter$count = 41797;
	#10 counter$count = 41798;
	#10 counter$count = 41799;
	#10 counter$count = 41800;
	#10 counter$count = 41801;
	#10 counter$count = 41802;
	#10 counter$count = 41803;
	#10 counter$count = 41804;
	#10 counter$count = 41805;
	#10 counter$count = 41806;
	#10 counter$count = 41807;
	#10 counter$count = 41808;
	#10 counter$count = 41809;
	#10 counter$count = 41810;
	#10 counter$count = 41811;
	#10 counter$count = 41812;
	#10 counter$count = 41813;
	#10 counter$count = 41814;
	#10 counter$count = 41815;
	#10 counter$count = 41816;
	#10 counter$count = 41817;
	#10 counter$count = 41818;
	#10 counter$count = 41819;
	#10 counter$count = 41820;
	#10 counter$count = 41821;
	#10 counter$count = 41822;
	#10 counter$count = 41823;
	#10 counter$count = 41824;
	#10 counter$count = 41825;
	#10 counter$count = 41826;
	#10 counter$count = 41827;
	#10 counter$count = 41828;
	#10 counter$count = 41829;
	#10 counter$count = 41830;
	#10 counter$count = 41831;
	#10 counter$count = 41832;
	#10 counter$count = 41833;
	#10 counter$count = 41834;
	#10 counter$count = 41835;
	#10 counter$count = 41836;
	#10 counter$count = 41837;
	#10 counter$count = 41838;
	#10 counter$count = 41839;
	#10 counter$count = 41840;
	#10 counter$count = 41841;
	#10 counter$count = 41842;
	#10 counter$count = 41843;
	#10 counter$count = 41844;
	#10 counter$count = 41845;
	#10 counter$count = 41846;
	#10 counter$count = 41847;
	#10 counter$count = 41848;
	#10 counter$count = 41849;
	#10 counter$count = 41850;
	#10 counter$count = 41851;
	#10 counter$count = 41852;
	#10 counter$count = 41853;
	#10 counter$count = 41854;
	#10 counter$count = 41855;
	#10 counter$count = 41856;
	#10 counter$count = 41857;
	#10 counter$count = 41858;
	#10 counter$count = 41859;
	#10 counter$count = 41860;
	#10 counter$count = 41861;
	#10 counter$count = 41862;
	#10 counter$count = 41863;
	#10 counter$count = 41864;
	#10 counter$count = 41865;
	#10 counter$count = 41866;
	#10 counter$count = 41867;
	#10 counter$count = 41868;
	#10 counter$count = 41869;
	#10 counter$count = 41870;
	#10 counter$count = 41871;
	#10 counter$count = 41872;
	#10 counter$count = 41873;
	#10 counter$count = 41874;
	#10 counter$count = 41875;
	#10 counter$count = 41876;
	#10 counter$count = 41877;
	#10 counter$count = 41878;
	#10 counter$count = 41879;
	#10 counter$count = 41880;
	#10 counter$count = 41881;
	#10 counter$count = 41882;
	#10 counter$count = 41883;
	#10 counter$count = 41884;
	#10 counter$count = 41885;
	#10 counter$count = 41886;
	#10 counter$count = 41887;
	#10 counter$count = 41888;
	#10 counter$count = 41889;
	#10 counter$count = 41890;
	#10 counter$count = 41891;
	#10 counter$count = 41892;
	#10 counter$count = 41893;
	#10 counter$count = 41894;
	#10 counter$count = 41895;
	#10 counter$count = 41896;
	#10 counter$count = 41897;
	#10 counter$count = 41898;
	#10 counter$count = 41899;
	#10 counter$count = 41900;
	#10 counter$count = 41901;
	#10 counter$count = 41902;
	#10 counter$count = 41903;
	#10 counter$count = 41904;
	#10 counter$count = 41905;
	#10 counter$count = 41906;
	#10 counter$count = 41907;
	#10 counter$count = 41908;
	#10 counter$count = 41909;
	#10 counter$count = 41910;
	#10 counter$count = 41911;
	#10 counter$count = 41912;
	#10 counter$count = 41913;
	#10 counter$count = 41914;
	#10 counter$count = 41915;
	#10 counter$count = 41916;
	#10 counter$count = 41917;
	#10 counter$count = 41918;
	#10 counter$count = 41919;
	#10 counter$count = 41920;
	#10 counter$count = 41921;
	#10 counter$count = 41922;
	#10 counter$count = 41923;
	#10 counter$count = 41924;
	#10 counter$count = 41925;
	#10 counter$count = 41926;
	#10 counter$count = 41927;
	#10 counter$count = 41928;
	#10 counter$count = 41929;
	#10 counter$count = 41930;
	#10 counter$count = 41931;
	#10 counter$count = 41932;
	#10 counter$count = 41933;
	#10 counter$count = 41934;
	#10 counter$count = 41935;
	#10 counter$count = 41936;
	#10 counter$count = 41937;
	#10 counter$count = 41938;
	#10 counter$count = 41939;
	#10 counter$count = 41940;
	#10 counter$count = 41941;
	#10 counter$count = 41942;
	#10 counter$count = 41943;
	#10 counter$count = 41944;
	#10 counter$count = 41945;
	#10 counter$count = 41946;
	#10 counter$count = 41947;
	#10 counter$count = 41948;
	#10 counter$count = 41949;
	#10 counter$count = 41950;
	#10 counter$count = 41951;
	#10 counter$count = 41952;
	#10 counter$count = 41953;
	#10 counter$count = 41954;
	#10 counter$count = 41955;
	#10 counter$count = 41956;
	#10 counter$count = 41957;
	#10 counter$count = 41958;
	#10 counter$count = 41959;
	#10 counter$count = 41960;
	#10 counter$count = 41961;
	#10 counter$count = 41962;
	#10 counter$count = 41963;
	#10 counter$count = 41964;
	#10 counter$count = 41965;
	#10 counter$count = 41966;
	#10 counter$count = 41967;
	#10 counter$count = 41968;
	#10 counter$count = 41969;
	#10 counter$count = 41970;
	#10 counter$count = 41971;
	#10 counter$count = 41972;
	#10 counter$count = 41973;
	#10 counter$count = 41974;
	#10 counter$count = 41975;
	#10 counter$count = 41976;
	#10 counter$count = 41977;
	#10 counter$count = 41978;
	#10 counter$count = 41979;
	#10 counter$count = 41980;
	#10 counter$count = 41981;
	#10 counter$count = 41982;
	#10 counter$count = 41983;
	#10 counter$count = 41984;
	#10 counter$count = 41985;
	#10 counter$count = 41986;
	#10 counter$count = 41987;
	#10 counter$count = 41988;
	#10 counter$count = 41989;
	#10 counter$count = 41990;
	#10 counter$count = 41991;
	#10 counter$count = 41992;
	#10 counter$count = 41993;
	#10 counter$count = 41994;
	#10 counter$count = 41995;
	#10 counter$count = 41996;
	#10 counter$count = 41997;
	#10 counter$count = 41998;
	#10 counter$count = 41999;
	#10 counter$count = 42000;
	#10 counter$count = 42001;
	#10 counter$count = 42002;
	#10 counter$count = 42003;
	#10 counter$count = 42004;
	#10 counter$count = 42005;
	#10 counter$count = 42006;
	#10 counter$count = 42007;
	#10 counter$count = 42008;
	#10 counter$count = 42009;
	#10 counter$count = 42010;
	#10 counter$count = 42011;
	#10 counter$count = 42012;
	#10 counter$count = 42013;
	#10 counter$count = 42014;
	#10 counter$count = 42015;
	#10 counter$count = 42016;
	#10 counter$count = 42017;
	#10 counter$count = 42018;
	#10 counter$count = 42019;
	#10 counter$count = 42020;
	#10 counter$count = 42021;
	#10 counter$count = 42022;
	#10 counter$count = 42023;
	#10 counter$count = 42024;
	#10 counter$count = 42025;
	#10 counter$count = 42026;
	#10 counter$count = 42027;
	#10 counter$count = 42028;
	#10 counter$count = 42029;
	#10 counter$count = 42030;
	#10 counter$count = 42031;
	#10 counter$count = 42032;
	#10 counter$count = 42033;
	#10 counter$count = 42034;
	#10 counter$count = 42035;
	#10 counter$count = 42036;
	#10 counter$count = 42037;
	#10 counter$count = 42038;
	#10 counter$count = 42039;
	#10 counter$count = 42040;
	#10 counter$count = 42041;
	#10 counter$count = 42042;
	#10 counter$count = 42043;
	#10 counter$count = 42044;
	#10 counter$count = 42045;
	#10 counter$count = 42046;
	#10 counter$count = 42047;
	#10 counter$count = 42048;
	#10 counter$count = 42049;
	#10 counter$count = 42050;
	#10 counter$count = 42051;
	#10 counter$count = 42052;
	#10 counter$count = 42053;
	#10 counter$count = 42054;
	#10 counter$count = 42055;
	#10 counter$count = 42056;
	#10 counter$count = 42057;
	#10 counter$count = 42058;
	#10 counter$count = 42059;
	#10 counter$count = 42060;
	#10 counter$count = 42061;
	#10 counter$count = 42062;
	#10 counter$count = 42063;
	#10 counter$count = 42064;
	#10 counter$count = 42065;
	#10 counter$count = 42066;
	#10 counter$count = 42067;
	#10 counter$count = 42068;
	#10 counter$count = 42069;
	#10 counter$count = 42070;
	#10 counter$count = 42071;
	#10 counter$count = 42072;
	#10 counter$count = 42073;
	#10 counter$count = 42074;
	#10 counter$count = 42075;
	#10 counter$count = 42076;
	#10 counter$count = 42077;
	#10 counter$count = 42078;
	#10 counter$count = 42079;
	#10 counter$count = 42080;
	#10 counter$count = 42081;
	#10 counter$count = 42082;
	#10 counter$count = 42083;
	#10 counter$count = 42084;
	#10 counter$count = 42085;
	#10 counter$count = 42086;
	#10 counter$count = 42087;
	#10 counter$count = 42088;
	#10 counter$count = 42089;
	#10 counter$count = 42090;
	#10 counter$count = 42091;
	#10 counter$count = 42092;
	#10 counter$count = 42093;
	#10 counter$count = 42094;
	#10 counter$count = 42095;
	#10 counter$count = 42096;
	#10 counter$count = 42097;
	#10 counter$count = 42098;
	#10 counter$count = 42099;
	#10 counter$count = 42100;
	#10 counter$count = 42101;
	#10 counter$count = 42102;
	#10 counter$count = 42103;
	#10 counter$count = 42104;
	#10 counter$count = 42105;
	#10 counter$count = 42106;
	#10 counter$count = 42107;
	#10 counter$count = 42108;
	#10 counter$count = 42109;
	#10 counter$count = 42110;
	#10 counter$count = 42111;
	#10 counter$count = 42112;
	#10 counter$count = 42113;
	#10 counter$count = 42114;
	#10 counter$count = 42115;
	#10 counter$count = 42116;
	#10 counter$count = 42117;
	#10 counter$count = 42118;
	#10 counter$count = 42119;
	#10 counter$count = 42120;
	#10 counter$count = 42121;
	#10 counter$count = 42122;
	#10 counter$count = 42123;
	#10 counter$count = 42124;
	#10 counter$count = 42125;
	#10 counter$count = 42126;
	#10 counter$count = 42127;
	#10 counter$count = 42128;
	#10 counter$count = 42129;
	#10 counter$count = 42130;
	#10 counter$count = 42131;
	#10 counter$count = 42132;
	#10 counter$count = 42133;
	#10 counter$count = 42134;
	#10 counter$count = 42135;
	#10 counter$count = 42136;
	#10 counter$count = 42137;
	#10 counter$count = 42138;
	#10 counter$count = 42139;
	#10 counter$count = 42140;
	#10 counter$count = 42141;
	#10 counter$count = 42142;
	#10 counter$count = 42143;
	#10 counter$count = 42144;
	#10 counter$count = 42145;
	#10 counter$count = 42146;
	#10 counter$count = 42147;
	#10 counter$count = 42148;
	#10 counter$count = 42149;
	#10 counter$count = 42150;
	#10 counter$count = 42151;
	#10 counter$count = 42152;
	#10 counter$count = 42153;
	#10 counter$count = 42154;
	#10 counter$count = 42155;
	#10 counter$count = 42156;
	#10 counter$count = 42157;
	#10 counter$count = 42158;
	#10 counter$count = 42159;
	#10 counter$count = 42160;
	#10 counter$count = 42161;
	#10 counter$count = 42162;
	#10 counter$count = 42163;
	#10 counter$count = 42164;
	#10 counter$count = 42165;
	#10 counter$count = 42166;
	#10 counter$count = 42167;
	#10 counter$count = 42168;
	#10 counter$count = 42169;
	#10 counter$count = 42170;
	#10 counter$count = 42171;
	#10 counter$count = 42172;
	#10 counter$count = 42173;
	#10 counter$count = 42174;
	#10 counter$count = 42175;
	#10 counter$count = 42176;
	#10 counter$count = 42177;
	#10 counter$count = 42178;
	#10 counter$count = 42179;
	#10 counter$count = 42180;
	#10 counter$count = 42181;
	#10 counter$count = 42182;
	#10 counter$count = 42183;
	#10 counter$count = 42184;
	#10 counter$count = 42185;
	#10 counter$count = 42186;
	#10 counter$count = 42187;
	#10 counter$count = 42188;
	#10 counter$count = 42189;
	#10 counter$count = 42190;
	#10 counter$count = 42191;
	#10 counter$count = 42192;
	#10 counter$count = 42193;
	#10 counter$count = 42194;
	#10 counter$count = 42195;
	#10 counter$count = 42196;
	#10 counter$count = 42197;
	#10 counter$count = 42198;
	#10 counter$count = 42199;
	#10 counter$count = 42200;
	#10 counter$count = 42201;
	#10 counter$count = 42202;
	#10 counter$count = 42203;
	#10 counter$count = 42204;
	#10 counter$count = 42205;
	#10 counter$count = 42206;
	#10 counter$count = 42207;
	#10 counter$count = 42208;
	#10 counter$count = 42209;
	#10 counter$count = 42210;
	#10 counter$count = 42211;
	#10 counter$count = 42212;
	#10 counter$count = 42213;
	#10 counter$count = 42214;
	#10 counter$count = 42215;
	#10 counter$count = 42216;
	#10 counter$count = 42217;
	#10 counter$count = 42218;
	#10 counter$count = 42219;
	#10 counter$count = 42220;
	#10 counter$count = 42221;
	#10 counter$count = 42222;
	#10 counter$count = 42223;
	#10 counter$count = 42224;
	#10 counter$count = 42225;
	#10 counter$count = 42226;
	#10 counter$count = 42227;
	#10 counter$count = 42228;
	#10 counter$count = 42229;
	#10 counter$count = 42230;
	#10 counter$count = 42231;
	#10 counter$count = 42232;
	#10 counter$count = 42233;
	#10 counter$count = 42234;
	#10 counter$count = 42235;
	#10 counter$count = 42236;
	#10 counter$count = 42237;
	#10 counter$count = 42238;
	#10 counter$count = 42239;
	#10 counter$count = 42240;
	#10 counter$count = 42241;
	#10 counter$count = 42242;
	#10 counter$count = 42243;
	#10 counter$count = 42244;
	#10 counter$count = 42245;
	#10 counter$count = 42246;
	#10 counter$count = 42247;
	#10 counter$count = 42248;
	#10 counter$count = 42249;
	#10 counter$count = 42250;
	#10 counter$count = 42251;
	#10 counter$count = 42252;
	#10 counter$count = 42253;
	#10 counter$count = 42254;
	#10 counter$count = 42255;
	#10 counter$count = 42256;
	#10 counter$count = 42257;
	#10 counter$count = 42258;
	#10 counter$count = 42259;
	#10 counter$count = 42260;
	#10 counter$count = 42261;
	#10 counter$count = 42262;
	#10 counter$count = 42263;
	#10 counter$count = 42264;
	#10 counter$count = 42265;
	#10 counter$count = 42266;
	#10 counter$count = 42267;
	#10 counter$count = 42268;
	#10 counter$count = 42269;
	#10 counter$count = 42270;
	#10 counter$count = 42271;
	#10 counter$count = 42272;
	#10 counter$count = 42273;
	#10 counter$count = 42274;
	#10 counter$count = 42275;
	#10 counter$count = 42276;
	#10 counter$count = 42277;
	#10 counter$count = 42278;
	#10 counter$count = 42279;
	#10 counter$count = 42280;
	#10 counter$count = 42281;
	#10 counter$count = 42282;
	#10 counter$count = 42283;
	#10 counter$count = 42284;
	#10 counter$count = 42285;
	#10 counter$count = 42286;
	#10 counter$count = 42287;
	#10 counter$count = 42288;
	#10 counter$count = 42289;
	#10 counter$count = 42290;
	#10 counter$count = 42291;
	#10 counter$count = 42292;
	#10 counter$count = 42293;
	#10 counter$count = 42294;
	#10 counter$count = 42295;
	#10 counter$count = 42296;
	#10 counter$count = 42297;
	#10 counter$count = 42298;
	#10 counter$count = 42299;
	#10 counter$count = 42300;
	#10 counter$count = 42301;
	#10 counter$count = 42302;
	#10 counter$count = 42303;
	#10 counter$count = 42304;
	#10 counter$count = 42305;
	#10 counter$count = 42306;
	#10 counter$count = 42307;
	#10 counter$count = 42308;
	#10 counter$count = 42309;
	#10 counter$count = 42310;
	#10 counter$count = 42311;
	#10 counter$count = 42312;
	#10 counter$count = 42313;
	#10 counter$count = 42314;
	#10 counter$count = 42315;
	#10 counter$count = 42316;
	#10 counter$count = 42317;
	#10 counter$count = 42318;
	#10 counter$count = 42319;
	#10 counter$count = 42320;
	#10 counter$count = 42321;
	#10 counter$count = 42322;
	#10 counter$count = 42323;
	#10 counter$count = 42324;
	#10 counter$count = 42325;
	#10 counter$count = 42326;
	#10 counter$count = 42327;
	#10 counter$count = 42328;
	#10 counter$count = 42329;
	#10 counter$count = 42330;
	#10 counter$count = 42331;
	#10 counter$count = 42332;
	#10 counter$count = 42333;
	#10 counter$count = 42334;
	#10 counter$count = 42335;
	#10 counter$count = 42336;
	#10 counter$count = 42337;
	#10 counter$count = 42338;
	#10 counter$count = 42339;
	#10 counter$count = 42340;
	#10 counter$count = 42341;
	#10 counter$count = 42342;
	#10 counter$count = 42343;
	#10 counter$count = 42344;
	#10 counter$count = 42345;
	#10 counter$count = 42346;
	#10 counter$count = 42347;
	#10 counter$count = 42348;
	#10 counter$count = 42349;
	#10 counter$count = 42350;
	#10 counter$count = 42351;
	#10 counter$count = 42352;
	#10 counter$count = 42353;
	#10 counter$count = 42354;
	#10 counter$count = 42355;
	#10 counter$count = 42356;
	#10 counter$count = 42357;
	#10 counter$count = 42358;
	#10 counter$count = 42359;
	#10 counter$count = 42360;
	#10 counter$count = 42361;
	#10 counter$count = 42362;
	#10 counter$count = 42363;
	#10 counter$count = 42364;
	#10 counter$count = 42365;
	#10 counter$count = 42366;
	#10 counter$count = 42367;
	#10 counter$count = 42368;
	#10 counter$count = 42369;
	#10 counter$count = 42370;
	#10 counter$count = 42371;
	#10 counter$count = 42372;
	#10 counter$count = 42373;
	#10 counter$count = 42374;
	#10 counter$count = 42375;
	#10 counter$count = 42376;
	#10 counter$count = 42377;
	#10 counter$count = 42378;
	#10 counter$count = 42379;
	#10 counter$count = 42380;
	#10 counter$count = 42381;
	#10 counter$count = 42382;
	#10 counter$count = 42383;
	#10 counter$count = 42384;
	#10 counter$count = 42385;
	#10 counter$count = 42386;
	#10 counter$count = 42387;
	#10 counter$count = 42388;
	#10 counter$count = 42389;
	#10 counter$count = 42390;
	#10 counter$count = 42391;
	#10 counter$count = 42392;
	#10 counter$count = 42393;
	#10 counter$count = 42394;
	#10 counter$count = 42395;
	#10 counter$count = 42396;
	#10 counter$count = 42397;
	#10 counter$count = 42398;
	#10 counter$count = 42399;
	#10 counter$count = 42400;
	#10 counter$count = 42401;
	#10 counter$count = 42402;
	#10 counter$count = 42403;
	#10 counter$count = 42404;
	#10 counter$count = 42405;
	#10 counter$count = 42406;
	#10 counter$count = 42407;
	#10 counter$count = 42408;
	#10 counter$count = 42409;
	#10 counter$count = 42410;
	#10 counter$count = 42411;
	#10 counter$count = 42412;
	#10 counter$count = 42413;
	#10 counter$count = 42414;
	#10 counter$count = 42415;
	#10 counter$count = 42416;
	#10 counter$count = 42417;
	#10 counter$count = 42418;
	#10 counter$count = 42419;
	#10 counter$count = 42420;
	#10 counter$count = 42421;
	#10 counter$count = 42422;
	#10 counter$count = 42423;
	#10 counter$count = 42424;
	#10 counter$count = 42425;
	#10 counter$count = 42426;
	#10 counter$count = 42427;
	#10 counter$count = 42428;
	#10 counter$count = 42429;
	#10 counter$count = 42430;
	#10 counter$count = 42431;
	#10 counter$count = 42432;
	#10 counter$count = 42433;
	#10 counter$count = 42434;
	#10 counter$count = 42435;
	#10 counter$count = 42436;
	#10 counter$count = 42437;
	#10 counter$count = 42438;
	#10 counter$count = 42439;
	#10 counter$count = 42440;
	#10 counter$count = 42441;
	#10 counter$count = 42442;
	#10 counter$count = 42443;
	#10 counter$count = 42444;
	#10 counter$count = 42445;
	#10 counter$count = 42446;
	#10 counter$count = 42447;
	#10 counter$count = 42448;
	#10 counter$count = 42449;
	#10 counter$count = 42450;
	#10 counter$count = 42451;
	#10 counter$count = 42452;
	#10 counter$count = 42453;
	#10 counter$count = 42454;
	#10 counter$count = 42455;
	#10 counter$count = 42456;
	#10 counter$count = 42457;
	#10 counter$count = 42458;
	#10 counter$count = 42459;
	#10 counter$count = 42460;
	#10 counter$count = 42461;
	#10 counter$count = 42462;
	#10 counter$count = 42463;
	#10 counter$count = 42464;
	#10 counter$count = 42465;
	#10 counter$count = 42466;
	#10 counter$count = 42467;
	#10 counter$count = 42468;
	#10 counter$count = 42469;
	#10 counter$count = 42470;
	#10 counter$count = 42471;
	#10 counter$count = 42472;
	#10 counter$count = 42473;
	#10 counter$count = 42474;
	#10 counter$count = 42475;
	#10 counter$count = 42476;
	#10 counter$count = 42477;
	#10 counter$count = 42478;
	#10 counter$count = 42479;
	#10 counter$count = 42480;
	#10 counter$count = 42481;
	#10 counter$count = 42482;
	#10 counter$count = 42483;
	#10 counter$count = 42484;
	#10 counter$count = 42485;
	#10 counter$count = 42486;
	#10 counter$count = 42487;
	#10 counter$count = 42488;
	#10 counter$count = 42489;
	#10 counter$count = 42490;
	#10 counter$count = 42491;
	#10 counter$count = 42492;
	#10 counter$count = 42493;
	#10 counter$count = 42494;
	#10 counter$count = 42495;
	#10 counter$count = 42496;
	#10 counter$count = 42497;
	#10 counter$count = 42498;
	#10 counter$count = 42499;
	#10 counter$count = 42500;
	#10 counter$count = 42501;
	#10 counter$count = 42502;
	#10 counter$count = 42503;
	#10 counter$count = 42504;
	#10 counter$count = 42505;
	#10 counter$count = 42506;
	#10 counter$count = 42507;
	#10 counter$count = 42508;
	#10 counter$count = 42509;
	#10 counter$count = 42510;
	#10 counter$count = 42511;
	#10 counter$count = 42512;
	#10 counter$count = 42513;
	#10 counter$count = 42514;
	#10 counter$count = 42515;
	#10 counter$count = 42516;
	#10 counter$count = 42517;
	#10 counter$count = 42518;
	#10 counter$count = 42519;
	#10 counter$count = 42520;
	#10 counter$count = 42521;
	#10 counter$count = 42522;
	#10 counter$count = 42523;
	#10 counter$count = 42524;
	#10 counter$count = 42525;
	#10 counter$count = 42526;
	#10 counter$count = 42527;
	#10 counter$count = 42528;
	#10 counter$count = 42529;
	#10 counter$count = 42530;
	#10 counter$count = 42531;
	#10 counter$count = 42532;
	#10 counter$count = 42533;
	#10 counter$count = 42534;
	#10 counter$count = 42535;
	#10 counter$count = 42536;
	#10 counter$count = 42537;
	#10 counter$count = 42538;
	#10 counter$count = 42539;
	#10 counter$count = 42540;
	#10 counter$count = 42541;
	#10 counter$count = 42542;
	#10 counter$count = 42543;
	#10 counter$count = 42544;
	#10 counter$count = 42545;
	#10 counter$count = 42546;
	#10 counter$count = 42547;
	#10 counter$count = 42548;
	#10 counter$count = 42549;
	#10 counter$count = 42550;
	#10 counter$count = 42551;
	#10 counter$count = 42552;
	#10 counter$count = 42553;
	#10 counter$count = 42554;
	#10 counter$count = 42555;
	#10 counter$count = 42556;
	#10 counter$count = 42557;
	#10 counter$count = 42558;
	#10 counter$count = 42559;
	#10 counter$count = 42560;
	#10 counter$count = 42561;
	#10 counter$count = 42562;
	#10 counter$count = 42563;
	#10 counter$count = 42564;
	#10 counter$count = 42565;
	#10 counter$count = 42566;
	#10 counter$count = 42567;
	#10 counter$count = 42568;
	#10 counter$count = 42569;
	#10 counter$count = 42570;
	#10 counter$count = 42571;
	#10 counter$count = 42572;
	#10 counter$count = 42573;
	#10 counter$count = 42574;
	#10 counter$count = 42575;
	#10 counter$count = 42576;
	#10 counter$count = 42577;
	#10 counter$count = 42578;
	#10 counter$count = 42579;
	#10 counter$count = 42580;
	#10 counter$count = 42581;
	#10 counter$count = 42582;
	#10 counter$count = 42583;
	#10 counter$count = 42584;
	#10 counter$count = 42585;
	#10 counter$count = 42586;
	#10 counter$count = 42587;
	#10 counter$count = 42588;
	#10 counter$count = 42589;
	#10 counter$count = 42590;
	#10 counter$count = 42591;
	#10 counter$count = 42592;
	#10 counter$count = 42593;
	#10 counter$count = 42594;
	#10 counter$count = 42595;
	#10 counter$count = 42596;
	#10 counter$count = 42597;
	#10 counter$count = 42598;
	#10 counter$count = 42599;
	#10 counter$count = 42600;
	#10 counter$count = 42601;
	#10 counter$count = 42602;
	#10 counter$count = 42603;
	#10 counter$count = 42604;
	#10 counter$count = 42605;
	#10 counter$count = 42606;
	#10 counter$count = 42607;
	#10 counter$count = 42608;
	#10 counter$count = 42609;
	#10 counter$count = 42610;
	#10 counter$count = 42611;
	#10 counter$count = 42612;
	#10 counter$count = 42613;
	#10 counter$count = 42614;
	#10 counter$count = 42615;
	#10 counter$count = 42616;
	#10 counter$count = 42617;
	#10 counter$count = 42618;
	#10 counter$count = 42619;
	#10 counter$count = 42620;
	#10 counter$count = 42621;
	#10 counter$count = 42622;
	#10 counter$count = 42623;
	#10 counter$count = 42624;
	#10 counter$count = 42625;
	#10 counter$count = 42626;
	#10 counter$count = 42627;
	#10 counter$count = 42628;
	#10 counter$count = 42629;
	#10 counter$count = 42630;
	#10 counter$count = 42631;
	#10 counter$count = 42632;
	#10 counter$count = 42633;
	#10 counter$count = 42634;
	#10 counter$count = 42635;
	#10 counter$count = 42636;
	#10 counter$count = 42637;
	#10 counter$count = 42638;
	#10 counter$count = 42639;
	#10 counter$count = 42640;
	#10 counter$count = 42641;
	#10 counter$count = 42642;
	#10 counter$count = 42643;
	#10 counter$count = 42644;
	#10 counter$count = 42645;
	#10 counter$count = 42646;
	#10 counter$count = 42647;
	#10 counter$count = 42648;
	#10 counter$count = 42649;
	#10 counter$count = 42650;
	#10 counter$count = 42651;
	#10 counter$count = 42652;
	#10 counter$count = 42653;
	#10 counter$count = 42654;
	#10 counter$count = 42655;
	#10 counter$count = 42656;
	#10 counter$count = 42657;
	#10 counter$count = 42658;
	#10 counter$count = 42659;
	#10 counter$count = 42660;
	#10 counter$count = 42661;
	#10 counter$count = 42662;
	#10 counter$count = 42663;
	#10 counter$count = 42664;
	#10 counter$count = 42665;
	#10 counter$count = 42666;
	#10 counter$count = 42667;
	#10 counter$count = 42668;
	#10 counter$count = 42669;
	#10 counter$count = 42670;
	#10 counter$count = 42671;
	#10 counter$count = 42672;
	#10 counter$count = 42673;
	#10 counter$count = 42674;
	#10 counter$count = 42675;
	#10 counter$count = 42676;
	#10 counter$count = 42677;
	#10 counter$count = 42678;
	#10 counter$count = 42679;
	#10 counter$count = 42680;
	#10 counter$count = 42681;
	#10 counter$count = 42682;
	#10 counter$count = 42683;
	#10 counter$count = 42684;
	#10 counter$count = 42685;
	#10 counter$count = 42686;
	#10 counter$count = 42687;
	#10 counter$count = 42688;
	#10 counter$count = 42689;
	#10 counter$count = 42690;
	#10 counter$count = 42691;
	#10 counter$count = 42692;
	#10 counter$count = 42693;
	#10 counter$count = 42694;
	#10 counter$count = 42695;
	#10 counter$count = 42696;
	#10 counter$count = 42697;
	#10 counter$count = 42698;
	#10 counter$count = 42699;
	#10 counter$count = 42700;
	#10 counter$count = 42701;
	#10 counter$count = 42702;
	#10 counter$count = 42703;
	#10 counter$count = 42704;
	#10 counter$count = 42705;
	#10 counter$count = 42706;
	#10 counter$count = 42707;
	#10 counter$count = 42708;
	#10 counter$count = 42709;
	#10 counter$count = 42710;
	#10 counter$count = 42711;
	#10 counter$count = 42712;
	#10 counter$count = 42713;
	#10 counter$count = 42714;
	#10 counter$count = 42715;
	#10 counter$count = 42716;
	#10 counter$count = 42717;
	#10 counter$count = 42718;
	#10 counter$count = 42719;
	#10 counter$count = 42720;
	#10 counter$count = 42721;
	#10 counter$count = 42722;
	#10 counter$count = 42723;
	#10 counter$count = 42724;
	#10 counter$count = 42725;
	#10 counter$count = 42726;
	#10 counter$count = 42727;
	#10 counter$count = 42728;
	#10 counter$count = 42729;
	#10 counter$count = 42730;
	#10 counter$count = 42731;
	#10 counter$count = 42732;
	#10 counter$count = 42733;
	#10 counter$count = 42734;
	#10 counter$count = 42735;
	#10 counter$count = 42736;
	#10 counter$count = 42737;
	#10 counter$count = 42738;
	#10 counter$count = 42739;
	#10 counter$count = 42740;
	#10 counter$count = 42741;
	#10 counter$count = 42742;
	#10 counter$count = 42743;
	#10 counter$count = 42744;
	#10 counter$count = 42745;
	#10 counter$count = 42746;
	#10 counter$count = 42747;
	#10 counter$count = 42748;
	#10 counter$count = 42749;
	#10 counter$count = 42750;
	#10 counter$count = 42751;
	#10 counter$count = 42752;
	#10 counter$count = 42753;
	#10 counter$count = 42754;
	#10 counter$count = 42755;
	#10 counter$count = 42756;
	#10 counter$count = 42757;
	#10 counter$count = 42758;
	#10 counter$count = 42759;
	#10 counter$count = 42760;
	#10 counter$count = 42761;
	#10 counter$count = 42762;
	#10 counter$count = 42763;
	#10 counter$count = 42764;
	#10 counter$count = 42765;
	#10 counter$count = 42766;
	#10 counter$count = 42767;
	#10 counter$count = 42768;
	#10 counter$count = 42769;
	#10 counter$count = 42770;
	#10 counter$count = 42771;
	#10 counter$count = 42772;
	#10 counter$count = 42773;
	#10 counter$count = 42774;
	#10 counter$count = 42775;
	#10 counter$count = 42776;
	#10 counter$count = 42777;
	#10 counter$count = 42778;
	#10 counter$count = 42779;
	#10 counter$count = 42780;
	#10 counter$count = 42781;
	#10 counter$count = 42782;
	#10 counter$count = 42783;
	#10 counter$count = 42784;
	#10 counter$count = 42785;
	#10 counter$count = 42786;
	#10 counter$count = 42787;
	#10 counter$count = 42788;
	#10 counter$count = 42789;
	#10 counter$count = 42790;
	#10 counter$count = 42791;
	#10 counter$count = 42792;
	#10 counter$count = 42793;
	#10 counter$count = 42794;
	#10 counter$count = 42795;
	#10 counter$count = 42796;
	#10 counter$count = 42797;
	#10 counter$count = 42798;
	#10 counter$count = 42799;
	#10 counter$count = 42800;
	#10 counter$count = 42801;
	#10 counter$count = 42802;
	#10 counter$count = 42803;
	#10 counter$count = 42804;
	#10 counter$count = 42805;
	#10 counter$count = 42806;
	#10 counter$count = 42807;
	#10 counter$count = 42808;
	#10 counter$count = 42809;
	#10 counter$count = 42810;
	#10 counter$count = 42811;
	#10 counter$count = 42812;
	#10 counter$count = 42813;
	#10 counter$count = 42814;
	#10 counter$count = 42815;
	#10 counter$count = 42816;
	#10 counter$count = 42817;
	#10 counter$count = 42818;
	#10 counter$count = 42819;
	#10 counter$count = 42820;
	#10 counter$count = 42821;
	#10 counter$count = 42822;
	#10 counter$count = 42823;
	#10 counter$count = 42824;
	#10 counter$count = 42825;
	#10 counter$count = 42826;
	#10 counter$count = 42827;
	#10 counter$count = 42828;
	#10 counter$count = 42829;
	#10 counter$count = 42830;
	#10 counter$count = 42831;
	#10 counter$count = 42832;
	#10 counter$count = 42833;
	#10 counter$count = 42834;
	#10 counter$count = 42835;
	#10 counter$count = 42836;
	#10 counter$count = 42837;
	#10 counter$count = 42838;
	#10 counter$count = 42839;
	#10 counter$count = 42840;
	#10 counter$count = 42841;
	#10 counter$count = 42842;
	#10 counter$count = 42843;
	#10 counter$count = 42844;
	#10 counter$count = 42845;
	#10 counter$count = 42846;
	#10 counter$count = 42847;
	#10 counter$count = 42848;
	#10 counter$count = 42849;
	#10 counter$count = 42850;
	#10 counter$count = 42851;
	#10 counter$count = 42852;
	#10 counter$count = 42853;
	#10 counter$count = 42854;
	#10 counter$count = 42855;
	#10 counter$count = 42856;
	#10 counter$count = 42857;
	#10 counter$count = 42858;
	#10 counter$count = 42859;
	#10 counter$count = 42860;
	#10 counter$count = 42861;
	#10 counter$count = 42862;
	#10 counter$count = 42863;
	#10 counter$count = 42864;
	#10 counter$count = 42865;
	#10 counter$count = 42866;
	#10 counter$count = 42867;
	#10 counter$count = 42868;
	#10 counter$count = 42869;
	#10 counter$count = 42870;
	#10 counter$count = 42871;
	#10 counter$count = 42872;
	#10 counter$count = 42873;
	#10 counter$count = 42874;
	#10 counter$count = 42875;
	#10 counter$count = 42876;
	#10 counter$count = 42877;
	#10 counter$count = 42878;
	#10 counter$count = 42879;
	#10 counter$count = 42880;
	#10 counter$count = 42881;
	#10 counter$count = 42882;
	#10 counter$count = 42883;
	#10 counter$count = 42884;
	#10 counter$count = 42885;
	#10 counter$count = 42886;
	#10 counter$count = 42887;
	#10 counter$count = 42888;
	#10 counter$count = 42889;
	#10 counter$count = 42890;
	#10 counter$count = 42891;
	#10 counter$count = 42892;
	#10 counter$count = 42893;
	#10 counter$count = 42894;
	#10 counter$count = 42895;
	#10 counter$count = 42896;
	#10 counter$count = 42897;
	#10 counter$count = 42898;
	#10 counter$count = 42899;
	#10 counter$count = 42900;
	#10 counter$count = 42901;
	#10 counter$count = 42902;
	#10 counter$count = 42903;
	#10 counter$count = 42904;
	#10 counter$count = 42905;
	#10 counter$count = 42906;
	#10 counter$count = 42907;
	#10 counter$count = 42908;
	#10 counter$count = 42909;
	#10 counter$count = 42910;
	#10 counter$count = 42911;
	#10 counter$count = 42912;
	#10 counter$count = 42913;
	#10 counter$count = 42914;
	#10 counter$count = 42915;
	#10 counter$count = 42916;
	#10 counter$count = 42917;
	#10 counter$count = 42918;
	#10 counter$count = 42919;
	#10 counter$count = 42920;
	#10 counter$count = 42921;
	#10 counter$count = 42922;
	#10 counter$count = 42923;
	#10 counter$count = 42924;
	#10 counter$count = 42925;
	#10 counter$count = 42926;
	#10 counter$count = 42927;
	#10 counter$count = 42928;
	#10 counter$count = 42929;
	#10 counter$count = 42930;
	#10 counter$count = 42931;
	#10 counter$count = 42932;
	#10 counter$count = 42933;
	#10 counter$count = 42934;
	#10 counter$count = 42935;
	#10 counter$count = 42936;
	#10 counter$count = 42937;
	#10 counter$count = 42938;
	#10 counter$count = 42939;
	#10 counter$count = 42940;
	#10 counter$count = 42941;
	#10 counter$count = 42942;
	#10 counter$count = 42943;
	#10 counter$count = 42944;
	#10 counter$count = 42945;
	#10 counter$count = 42946;
	#10 counter$count = 42947;
	#10 counter$count = 42948;
	#10 counter$count = 42949;
	#10 counter$count = 42950;
	#10 counter$count = 42951;
	#10 counter$count = 42952;
	#10 counter$count = 42953;
	#10 counter$count = 42954;
	#10 counter$count = 42955;
	#10 counter$count = 42956;
	#10 counter$count = 42957;
	#10 counter$count = 42958;
	#10 counter$count = 42959;
	#10 counter$count = 42960;
	#10 counter$count = 42961;
	#10 counter$count = 42962;
	#10 counter$count = 42963;
	#10 counter$count = 42964;
	#10 counter$count = 42965;
	#10 counter$count = 42966;
	#10 counter$count = 42967;
	#10 counter$count = 42968;
	#10 counter$count = 42969;
	#10 counter$count = 42970;
	#10 counter$count = 42971;
	#10 counter$count = 42972;
	#10 counter$count = 42973;
	#10 counter$count = 42974;
	#10 counter$count = 42975;
	#10 counter$count = 42976;
	#10 counter$count = 42977;
	#10 counter$count = 42978;
	#10 counter$count = 42979;
	#10 counter$count = 42980;
	#10 counter$count = 42981;
	#10 counter$count = 42982;
	#10 counter$count = 42983;
	#10 counter$count = 42984;
	#10 counter$count = 42985;
	#10 counter$count = 42986;
	#10 counter$count = 42987;
	#10 counter$count = 42988;
	#10 counter$count = 42989;
	#10 counter$count = 42990;
	#10 counter$count = 42991;
	#10 counter$count = 42992;
	#10 counter$count = 42993;
	#10 counter$count = 42994;
	#10 counter$count = 42995;
	#10 counter$count = 42996;
	#10 counter$count = 42997;
	#10 counter$count = 42998;
	#10 counter$count = 42999;
	#10 counter$count = 43000;
	#10 counter$count = 43001;
	#10 counter$count = 43002;
	#10 counter$count = 43003;
	#10 counter$count = 43004;
	#10 counter$count = 43005;
	#10 counter$count = 43006;
	#10 counter$count = 43007;
	#10 counter$count = 43008;
	#10 counter$count = 43009;
	#10 counter$count = 43010;
	#10 counter$count = 43011;
	#10 counter$count = 43012;
	#10 counter$count = 43013;
	#10 counter$count = 43014;
	#10 counter$count = 43015;
	#10 counter$count = 43016;
	#10 counter$count = 43017;
	#10 counter$count = 43018;
	#10 counter$count = 43019;
	#10 counter$count = 43020;
	#10 counter$count = 43021;
	#10 counter$count = 43022;
	#10 counter$count = 43023;
	#10 counter$count = 43024;
	#10 counter$count = 43025;
	#10 counter$count = 43026;
	#10 counter$count = 43027;
	#10 counter$count = 43028;
	#10 counter$count = 43029;
	#10 counter$count = 43030;
	#10 counter$count = 43031;
	#10 counter$count = 43032;
	#10 counter$count = 43033;
	#10 counter$count = 43034;
	#10 counter$count = 43035;
	#10 counter$count = 43036;
	#10 counter$count = 43037;
	#10 counter$count = 43038;
	#10 counter$count = 43039;
	#10 counter$count = 43040;
	#10 counter$count = 43041;
	#10 counter$count = 43042;
	#10 counter$count = 43043;
	#10 counter$count = 43044;
	#10 counter$count = 43045;
	#10 counter$count = 43046;
	#10 counter$count = 43047;
	#10 counter$count = 43048;
	#10 counter$count = 43049;
	#10 counter$count = 43050;
	#10 counter$count = 43051;
	#10 counter$count = 43052;
	#10 counter$count = 43053;
	#10 counter$count = 43054;
	#10 counter$count = 43055;
	#10 counter$count = 43056;
	#10 counter$count = 43057;
	#10 counter$count = 43058;
	#10 counter$count = 43059;
	#10 counter$count = 43060;
	#10 counter$count = 43061;
	#10 counter$count = 43062;
	#10 counter$count = 43063;
	#10 counter$count = 43064;
	#10 counter$count = 43065;
	#10 counter$count = 43066;
	#10 counter$count = 43067;
	#10 counter$count = 43068;
	#10 counter$count = 43069;
	#10 counter$count = 43070;
	#10 counter$count = 43071;
	#10 counter$count = 43072;
	#10 counter$count = 43073;
	#10 counter$count = 43074;
	#10 counter$count = 43075;
	#10 counter$count = 43076;
	#10 counter$count = 43077;
	#10 counter$count = 43078;
	#10 counter$count = 43079;
	#10 counter$count = 43080;
	#10 counter$count = 43081;
	#10 counter$count = 43082;
	#10 counter$count = 43083;
	#10 counter$count = 43084;
	#10 counter$count = 43085;
	#10 counter$count = 43086;
	#10 counter$count = 43087;
	#10 counter$count = 43088;
	#10 counter$count = 43089;
	#10 counter$count = 43090;
	#10 counter$count = 43091;
	#10 counter$count = 43092;
	#10 counter$count = 43093;
	#10 counter$count = 43094;
	#10 counter$count = 43095;
	#10 counter$count = 43096;
	#10 counter$count = 43097;
	#10 counter$count = 43098;
	#10 counter$count = 43099;
	#10 counter$count = 43100;
	#10 counter$count = 43101;
	#10 counter$count = 43102;
	#10 counter$count = 43103;
	#10 counter$count = 43104;
	#10 counter$count = 43105;
	#10 counter$count = 43106;
	#10 counter$count = 43107;
	#10 counter$count = 43108;
	#10 counter$count = 43109;
	#10 counter$count = 43110;
	#10 counter$count = 43111;
	#10 counter$count = 43112;
	#10 counter$count = 43113;
	#10 counter$count = 43114;
	#10 counter$count = 43115;
	#10 counter$count = 43116;
	#10 counter$count = 43117;
	#10 counter$count = 43118;
	#10 counter$count = 43119;
	#10 counter$count = 43120;
	#10 counter$count = 43121;
	#10 counter$count = 43122;
	#10 counter$count = 43123;
	#10 counter$count = 43124;
	#10 counter$count = 43125;
	#10 counter$count = 43126;
	#10 counter$count = 43127;
	#10 counter$count = 43128;
	#10 counter$count = 43129;
	#10 counter$count = 43130;
	#10 counter$count = 43131;
	#10 counter$count = 43132;
	#10 counter$count = 43133;
	#10 counter$count = 43134;
	#10 counter$count = 43135;
	#10 counter$count = 43136;
	#10 counter$count = 43137;
	#10 counter$count = 43138;
	#10 counter$count = 43139;
	#10 counter$count = 43140;
	#10 counter$count = 43141;
	#10 counter$count = 43142;
	#10 counter$count = 43143;
	#10 counter$count = 43144;
	#10 counter$count = 43145;
	#10 counter$count = 43146;
	#10 counter$count = 43147;
	#10 counter$count = 43148;
	#10 counter$count = 43149;
	#10 counter$count = 43150;
	#10 counter$count = 43151;
	#10 counter$count = 43152;
	#10 counter$count = 43153;
	#10 counter$count = 43154;
	#10 counter$count = 43155;
	#10 counter$count = 43156;
	#10 counter$count = 43157;
	#10 counter$count = 43158;
	#10 counter$count = 43159;
	#10 counter$count = 43160;
	#10 counter$count = 43161;
	#10 counter$count = 43162;
	#10 counter$count = 43163;
	#10 counter$count = 43164;
	#10 counter$count = 43165;
	#10 counter$count = 43166;
	#10 counter$count = 43167;
	#10 counter$count = 43168;
	#10 counter$count = 43169;
	#10 counter$count = 43170;
	#10 counter$count = 43171;
	#10 counter$count = 43172;
	#10 counter$count = 43173;
	#10 counter$count = 43174;
	#10 counter$count = 43175;
	#10 counter$count = 43176;
	#10 counter$count = 43177;
	#10 counter$count = 43178;
	#10 counter$count = 43179;
	#10 counter$count = 43180;
	#10 counter$count = 43181;
	#10 counter$count = 43182;
	#10 counter$count = 43183;
	#10 counter$count = 43184;
	#10 counter$count = 43185;
	#10 counter$count = 43186;
	#10 counter$count = 43187;
	#10 counter$count = 43188;
	#10 counter$count = 43189;
	#10 counter$count = 43190;
	#10 counter$count = 43191;
	#10 counter$count = 43192;
	#10 counter$count = 43193;
	#10 counter$count = 43194;
	#10 counter$count = 43195;
	#10 counter$count = 43196;
	#10 counter$count = 43197;
	#10 counter$count = 43198;
	#10 counter$count = 43199;
	#10 counter$count = 43200;
	#10 counter$count = 43201;
	#10 counter$count = 43202;
	#10 counter$count = 43203;
	#10 counter$count = 43204;
	#10 counter$count = 43205;
	#10 counter$count = 43206;
	#10 counter$count = 43207;
	#10 counter$count = 43208;
	#10 counter$count = 43209;
	#10 counter$count = 43210;
	#10 counter$count = 43211;
	#10 counter$count = 43212;
	#10 counter$count = 43213;
	#10 counter$count = 43214;
	#10 counter$count = 43215;
	#10 counter$count = 43216;
	#10 counter$count = 43217;
	#10 counter$count = 43218;
	#10 counter$count = 43219;
	#10 counter$count = 43220;
	#10 counter$count = 43221;
	#10 counter$count = 43222;
	#10 counter$count = 43223;
	#10 counter$count = 43224;
	#10 counter$count = 43225;
	#10 counter$count = 43226;
	#10 counter$count = 43227;
	#10 counter$count = 43228;
	#10 counter$count = 43229;
	#10 counter$count = 43230;
	#10 counter$count = 43231;
	#10 counter$count = 43232;
	#10 counter$count = 43233;
	#10 counter$count = 43234;
	#10 counter$count = 43235;
	#10 counter$count = 43236;
	#10 counter$count = 43237;
	#10 counter$count = 43238;
	#10 counter$count = 43239;
	#10 counter$count = 43240;
	#10 counter$count = 43241;
	#10 counter$count = 43242;
	#10 counter$count = 43243;
	#10 counter$count = 43244;
	#10 counter$count = 43245;
	#10 counter$count = 43246;
	#10 counter$count = 43247;
	#10 counter$count = 43248;
	#10 counter$count = 43249;
	#10 counter$count = 43250;
	#10 counter$count = 43251;
	#10 counter$count = 43252;
	#10 counter$count = 43253;
	#10 counter$count = 43254;
	#10 counter$count = 43255;
	#10 counter$count = 43256;
	#10 counter$count = 43257;
	#10 counter$count = 43258;
	#10 counter$count = 43259;
	#10 counter$count = 43260;
	#10 counter$count = 43261;
	#10 counter$count = 43262;
	#10 counter$count = 43263;
	#10 counter$count = 43264;
	#10 counter$count = 43265;
	#10 counter$count = 43266;
	#10 counter$count = 43267;
	#10 counter$count = 43268;
	#10 counter$count = 43269;
	#10 counter$count = 43270;
	#10 counter$count = 43271;
	#10 counter$count = 43272;
	#10 counter$count = 43273;
	#10 counter$count = 43274;
	#10 counter$count = 43275;
	#10 counter$count = 43276;
	#10 counter$count = 43277;
	#10 counter$count = 43278;
	#10 counter$count = 43279;
	#10 counter$count = 43280;
	#10 counter$count = 43281;
	#10 counter$count = 43282;
	#10 counter$count = 43283;
	#10 counter$count = 43284;
	#10 counter$count = 43285;
	#10 counter$count = 43286;
	#10 counter$count = 43287;
	#10 counter$count = 43288;
	#10 counter$count = 43289;
	#10 counter$count = 43290;
	#10 counter$count = 43291;
	#10 counter$count = 43292;
	#10 counter$count = 43293;
	#10 counter$count = 43294;
	#10 counter$count = 43295;
	#10 counter$count = 43296;
	#10 counter$count = 43297;
	#10 counter$count = 43298;
	#10 counter$count = 43299;
	#10 counter$count = 43300;
	#10 counter$count = 43301;
	#10 counter$count = 43302;
	#10 counter$count = 43303;
	#10 counter$count = 43304;
	#10 counter$count = 43305;
	#10 counter$count = 43306;
	#10 counter$count = 43307;
	#10 counter$count = 43308;
	#10 counter$count = 43309;
	#10 counter$count = 43310;
	#10 counter$count = 43311;
	#10 counter$count = 43312;
	#10 counter$count = 43313;
	#10 counter$count = 43314;
	#10 counter$count = 43315;
	#10 counter$count = 43316;
	#10 counter$count = 43317;
	#10 counter$count = 43318;
	#10 counter$count = 43319;
	#10 counter$count = 43320;
	#10 counter$count = 43321;
	#10 counter$count = 43322;
	#10 counter$count = 43323;
	#10 counter$count = 43324;
	#10 counter$count = 43325;
	#10 counter$count = 43326;
	#10 counter$count = 43327;
	#10 counter$count = 43328;
	#10 counter$count = 43329;
	#10 counter$count = 43330;
	#10 counter$count = 43331;
	#10 counter$count = 43332;
	#10 counter$count = 43333;
	#10 counter$count = 43334;
	#10 counter$count = 43335;
	#10 counter$count = 43336;
	#10 counter$count = 43337;
	#10 counter$count = 43338;
	#10 counter$count = 43339;
	#10 counter$count = 43340;
	#10 counter$count = 43341;
	#10 counter$count = 43342;
	#10 counter$count = 43343;
	#10 counter$count = 43344;
	#10 counter$count = 43345;
	#10 counter$count = 43346;
	#10 counter$count = 43347;
	#10 counter$count = 43348;
	#10 counter$count = 43349;
	#10 counter$count = 43350;
	#10 counter$count = 43351;
	#10 counter$count = 43352;
	#10 counter$count = 43353;
	#10 counter$count = 43354;
	#10 counter$count = 43355;
	#10 counter$count = 43356;
	#10 counter$count = 43357;
	#10 counter$count = 43358;
	#10 counter$count = 43359;
	#10 counter$count = 43360;
	#10 counter$count = 43361;
	#10 counter$count = 43362;
	#10 counter$count = 43363;
	#10 counter$count = 43364;
	#10 counter$count = 43365;
	#10 counter$count = 43366;
	#10 counter$count = 43367;
	#10 counter$count = 43368;
	#10 counter$count = 43369;
	#10 counter$count = 43370;
	#10 counter$count = 43371;
	#10 counter$count = 43372;
	#10 counter$count = 43373;
	#10 counter$count = 43374;
	#10 counter$count = 43375;
	#10 counter$count = 43376;
	#10 counter$count = 43377;
	#10 counter$count = 43378;
	#10 counter$count = 43379;
	#10 counter$count = 43380;
	#10 counter$count = 43381;
	#10 counter$count = 43382;
	#10 counter$count = 43383;
	#10 counter$count = 43384;
	#10 counter$count = 43385;
	#10 counter$count = 43386;
	#10 counter$count = 43387;
	#10 counter$count = 43388;
	#10 counter$count = 43389;
	#10 counter$count = 43390;
	#10 counter$count = 43391;
	#10 counter$count = 43392;
	#10 counter$count = 43393;
	#10 counter$count = 43394;
	#10 counter$count = 43395;
	#10 counter$count = 43396;
	#10 counter$count = 43397;
	#10 counter$count = 43398;
	#10 counter$count = 43399;
	#10 counter$count = 43400;
	#10 counter$count = 43401;
	#10 counter$count = 43402;
	#10 counter$count = 43403;
	#10 counter$count = 43404;
	#10 counter$count = 43405;
	#10 counter$count = 43406;
	#10 counter$count = 43407;
	#10 counter$count = 43408;
	#10 counter$count = 43409;
	#10 counter$count = 43410;
	#10 counter$count = 43411;
	#10 counter$count = 43412;
	#10 counter$count = 43413;
	#10 counter$count = 43414;
	#10 counter$count = 43415;
	#10 counter$count = 43416;
	#10 counter$count = 43417;
	#10 counter$count = 43418;
	#10 counter$count = 43419;
	#10 counter$count = 43420;
	#10 counter$count = 43421;
	#10 counter$count = 43422;
	#10 counter$count = 43423;
	#10 counter$count = 43424;
	#10 counter$count = 43425;
	#10 counter$count = 43426;
	#10 counter$count = 43427;
	#10 counter$count = 43428;
	#10 counter$count = 43429;
	#10 counter$count = 43430;
	#10 counter$count = 43431;
	#10 counter$count = 43432;
	#10 counter$count = 43433;
	#10 counter$count = 43434;
	#10 counter$count = 43435;
	#10 counter$count = 43436;
	#10 counter$count = 43437;
	#10 counter$count = 43438;
	#10 counter$count = 43439;
	#10 counter$count = 43440;
	#10 counter$count = 43441;
	#10 counter$count = 43442;
	#10 counter$count = 43443;
	#10 counter$count = 43444;
	#10 counter$count = 43445;
	#10 counter$count = 43446;
	#10 counter$count = 43447;
	#10 counter$count = 43448;
	#10 counter$count = 43449;
	#10 counter$count = 43450;
	#10 counter$count = 43451;
	#10 counter$count = 43452;
	#10 counter$count = 43453;
	#10 counter$count = 43454;
	#10 counter$count = 43455;
	#10 counter$count = 43456;
	#10 counter$count = 43457;
	#10 counter$count = 43458;
	#10 counter$count = 43459;
	#10 counter$count = 43460;
	#10 counter$count = 43461;
	#10 counter$count = 43462;
	#10 counter$count = 43463;
	#10 counter$count = 43464;
	#10 counter$count = 43465;
	#10 counter$count = 43466;
	#10 counter$count = 43467;
	#10 counter$count = 43468;
	#10 counter$count = 43469;
	#10 counter$count = 43470;
	#10 counter$count = 43471;
	#10 counter$count = 43472;
	#10 counter$count = 43473;
	#10 counter$count = 43474;
	#10 counter$count = 43475;
	#10 counter$count = 43476;
	#10 counter$count = 43477;
	#10 counter$count = 43478;
	#10 counter$count = 43479;
	#10 counter$count = 43480;
	#10 counter$count = 43481;
	#10 counter$count = 43482;
	#10 counter$count = 43483;
	#10 counter$count = 43484;
	#10 counter$count = 43485;
	#10 counter$count = 43486;
	#10 counter$count = 43487;
	#10 counter$count = 43488;
	#10 counter$count = 43489;
	#10 counter$count = 43490;
	#10 counter$count = 43491;
	#10 counter$count = 43492;
	#10 counter$count = 43493;
	#10 counter$count = 43494;
	#10 counter$count = 43495;
	#10 counter$count = 43496;
	#10 counter$count = 43497;
	#10 counter$count = 43498;
	#10 counter$count = 43499;
	#10 counter$count = 43500;
	#10 counter$count = 43501;
	#10 counter$count = 43502;
	#10 counter$count = 43503;
	#10 counter$count = 43504;
	#10 counter$count = 43505;
	#10 counter$count = 43506;
	#10 counter$count = 43507;
	#10 counter$count = 43508;
	#10 counter$count = 43509;
	#10 counter$count = 43510;
	#10 counter$count = 43511;
	#10 counter$count = 43512;
	#10 counter$count = 43513;
	#10 counter$count = 43514;
	#10 counter$count = 43515;
	#10 counter$count = 43516;
	#10 counter$count = 43517;
	#10 counter$count = 43518;
	#10 counter$count = 43519;
	#10 counter$count = 43520;
	#10 counter$count = 43521;
	#10 counter$count = 43522;
	#10 counter$count = 43523;
	#10 counter$count = 43524;
	#10 counter$count = 43525;
	#10 counter$count = 43526;
	#10 counter$count = 43527;
	#10 counter$count = 43528;
	#10 counter$count = 43529;
	#10 counter$count = 43530;
	#10 counter$count = 43531;
	#10 counter$count = 43532;
	#10 counter$count = 43533;
	#10 counter$count = 43534;
	#10 counter$count = 43535;
	#10 counter$count = 43536;
	#10 counter$count = 43537;
	#10 counter$count = 43538;
	#10 counter$count = 43539;
	#10 counter$count = 43540;
	#10 counter$count = 43541;
	#10 counter$count = 43542;
	#10 counter$count = 43543;
	#10 counter$count = 43544;
	#10 counter$count = 43545;
	#10 counter$count = 43546;
	#10 counter$count = 43547;
	#10 counter$count = 43548;
	#10 counter$count = 43549;
	#10 counter$count = 43550;
	#10 counter$count = 43551;
	#10 counter$count = 43552;
	#10 counter$count = 43553;
	#10 counter$count = 43554;
	#10 counter$count = 43555;
	#10 counter$count = 43556;
	#10 counter$count = 43557;
	#10 counter$count = 43558;
	#10 counter$count = 43559;
	#10 counter$count = 43560;
	#10 counter$count = 43561;
	#10 counter$count = 43562;
	#10 counter$count = 43563;
	#10 counter$count = 43564;
	#10 counter$count = 43565;
	#10 counter$count = 43566;
	#10 counter$count = 43567;
	#10 counter$count = 43568;
	#10 counter$count = 43569;
	#10 counter$count = 43570;
	#10 counter$count = 43571;
	#10 counter$count = 43572;
	#10 counter$count = 43573;
	#10 counter$count = 43574;
	#10 counter$count = 43575;
	#10 counter$count = 43576;
	#10 counter$count = 43577;
	#10 counter$count = 43578;
	#10 counter$count = 43579;
	#10 counter$count = 43580;
	#10 counter$count = 43581;
	#10 counter$count = 43582;
	#10 counter$count = 43583;
	#10 counter$count = 43584;
	#10 counter$count = 43585;
	#10 counter$count = 43586;
	#10 counter$count = 43587;
	#10 counter$count = 43588;
	#10 counter$count = 43589;
	#10 counter$count = 43590;
	#10 counter$count = 43591;
	#10 counter$count = 43592;
	#10 counter$count = 43593;
	#10 counter$count = 43594;
	#10 counter$count = 43595;
	#10 counter$count = 43596;
	#10 counter$count = 43597;
	#10 counter$count = 43598;
	#10 counter$count = 43599;
	#10 counter$count = 43600;
	#10 counter$count = 43601;
	#10 counter$count = 43602;
	#10 counter$count = 43603;
	#10 counter$count = 43604;
	#10 counter$count = 43605;
	#10 counter$count = 43606;
	#10 counter$count = 43607;
	#10 counter$count = 43608;
	#10 counter$count = 43609;
	#10 counter$count = 43610;
	#10 counter$count = 43611;
	#10 counter$count = 43612;
	#10 counter$count = 43613;
	#10 counter$count = 43614;
	#10 counter$count = 43615;
	#10 counter$count = 43616;
	#10 counter$count = 43617;
	#10 counter$count = 43618;
	#10 counter$count = 43619;
	#10 counter$count = 43620;
	#10 counter$count = 43621;
	#10 counter$count = 43622;
	#10 counter$count = 43623;
	#10 counter$count = 43624;
	#10 counter$count = 43625;
	#10 counter$count = 43626;
	#10 counter$count = 43627;
	#10 counter$count = 43628;
	#10 counter$count = 43629;
	#10 counter$count = 43630;
	#10 counter$count = 43631;
	#10 counter$count = 43632;
	#10 counter$count = 43633;
	#10 counter$count = 43634;
	#10 counter$count = 43635;
	#10 counter$count = 43636;
	#10 counter$count = 43637;
	#10 counter$count = 43638;
	#10 counter$count = 43639;
	#10 counter$count = 43640;
	#10 counter$count = 43641;
	#10 counter$count = 43642;
	#10 counter$count = 43643;
	#10 counter$count = 43644;
	#10 counter$count = 43645;
	#10 counter$count = 43646;
	#10 counter$count = 43647;
	#10 counter$count = 43648;
	#10 counter$count = 43649;
	#10 counter$count = 43650;
	#10 counter$count = 43651;
	#10 counter$count = 43652;
	#10 counter$count = 43653;
	#10 counter$count = 43654;
	#10 counter$count = 43655;
	#10 counter$count = 43656;
	#10 counter$count = 43657;
	#10 counter$count = 43658;
	#10 counter$count = 43659;
	#10 counter$count = 43660;
	#10 counter$count = 43661;
	#10 counter$count = 43662;
	#10 counter$count = 43663;
	#10 counter$count = 43664;
	#10 counter$count = 43665;
	#10 counter$count = 43666;
	#10 counter$count = 43667;
	#10 counter$count = 43668;
	#10 counter$count = 43669;
	#10 counter$count = 43670;
	#10 counter$count = 43671;
	#10 counter$count = 43672;
	#10 counter$count = 43673;
	#10 counter$count = 43674;
	#10 counter$count = 43675;
	#10 counter$count = 43676;
	#10 counter$count = 43677;
	#10 counter$count = 43678;
	#10 counter$count = 43679;
	#10 counter$count = 43680;
	#10 counter$count = 43681;
	#10 counter$count = 43682;
	#10 counter$count = 43683;
	#10 counter$count = 43684;
	#10 counter$count = 43685;
	#10 counter$count = 43686;
	#10 counter$count = 43687;
	#10 counter$count = 43688;
	#10 counter$count = 43689;
	#10 counter$count = 43690;
	#10 counter$count = 43691;
	#10 counter$count = 43692;
	#10 counter$count = 43693;
	#10 counter$count = 43694;
	#10 counter$count = 43695;
	#10 counter$count = 43696;
	#10 counter$count = 43697;
	#10 counter$count = 43698;
	#10 counter$count = 43699;
	#10 counter$count = 43700;
	#10 counter$count = 43701;
	#10 counter$count = 43702;
	#10 counter$count = 43703;
	#10 counter$count = 43704;
	#10 counter$count = 43705;
	#10 counter$count = 43706;
	#10 counter$count = 43707;
	#10 counter$count = 43708;
	#10 counter$count = 43709;
	#10 counter$count = 43710;
	#10 counter$count = 43711;
	#10 counter$count = 43712;
	#10 counter$count = 43713;
	#10 counter$count = 43714;
	#10 counter$count = 43715;
	#10 counter$count = 43716;
	#10 counter$count = 43717;
	#10 counter$count = 43718;
	#10 counter$count = 43719;
	#10 counter$count = 43720;
	#10 counter$count = 43721;
	#10 counter$count = 43722;
	#10 counter$count = 43723;
	#10 counter$count = 43724;
	#10 counter$count = 43725;
	#10 counter$count = 43726;
	#10 counter$count = 43727;
	#10 counter$count = 43728;
	#10 counter$count = 43729;
	#10 counter$count = 43730;
	#10 counter$count = 43731;
	#10 counter$count = 43732;
	#10 counter$count = 43733;
	#10 counter$count = 43734;
	#10 counter$count = 43735;
	#10 counter$count = 43736;
	#10 counter$count = 43737;
	#10 counter$count = 43738;
	#10 counter$count = 43739;
	#10 counter$count = 43740;
	#10 counter$count = 43741;
	#10 counter$count = 43742;
	#10 counter$count = 43743;
	#10 counter$count = 43744;
	#10 counter$count = 43745;
	#10 counter$count = 43746;
	#10 counter$count = 43747;
	#10 counter$count = 43748;
	#10 counter$count = 43749;
	#10 counter$count = 43750;
	#10 counter$count = 43751;
	#10 counter$count = 43752;
	#10 counter$count = 43753;
	#10 counter$count = 43754;
	#10 counter$count = 43755;
	#10 counter$count = 43756;
	#10 counter$count = 43757;
	#10 counter$count = 43758;
	#10 counter$count = 43759;
	#10 counter$count = 43760;
	#10 counter$count = 43761;
	#10 counter$count = 43762;
	#10 counter$count = 43763;
	#10 counter$count = 43764;
	#10 counter$count = 43765;
	#10 counter$count = 43766;
	#10 counter$count = 43767;
	#10 counter$count = 43768;
	#10 counter$count = 43769;
	#10 counter$count = 43770;
	#10 counter$count = 43771;
	#10 counter$count = 43772;
	#10 counter$count = 43773;
	#10 counter$count = 43774;
	#10 counter$count = 43775;
	#10 counter$count = 43776;
	#10 counter$count = 43777;
	#10 counter$count = 43778;
	#10 counter$count = 43779;
	#10 counter$count = 43780;
	#10 counter$count = 43781;
	#10 counter$count = 43782;
	#10 counter$count = 43783;
	#10 counter$count = 43784;
	#10 counter$count = 43785;
	#10 counter$count = 43786;
	#10 counter$count = 43787;
	#10 counter$count = 43788;
	#10 counter$count = 43789;
	#10 counter$count = 43790;
	#10 counter$count = 43791;
	#10 counter$count = 43792;
	#10 counter$count = 43793;
	#10 counter$count = 43794;
	#10 counter$count = 43795;
	#10 counter$count = 43796;
	#10 counter$count = 43797;
	#10 counter$count = 43798;
	#10 counter$count = 43799;
	#10 counter$count = 43800;
	#10 counter$count = 43801;
	#10 counter$count = 43802;
	#10 counter$count = 43803;
	#10 counter$count = 43804;
	#10 counter$count = 43805;
	#10 counter$count = 43806;
	#10 counter$count = 43807;
	#10 counter$count = 43808;
	#10 counter$count = 43809;
	#10 counter$count = 43810;
	#10 counter$count = 43811;
	#10 counter$count = 43812;
	#10 counter$count = 43813;
	#10 counter$count = 43814;
	#10 counter$count = 43815;
	#10 counter$count = 43816;
	#10 counter$count = 43817;
	#10 counter$count = 43818;
	#10 counter$count = 43819;
	#10 counter$count = 43820;
	#10 counter$count = 43821;
	#10 counter$count = 43822;
	#10 counter$count = 43823;
	#10 counter$count = 43824;
	#10 counter$count = 43825;
	#10 counter$count = 43826;
	#10 counter$count = 43827;
	#10 counter$count = 43828;
	#10 counter$count = 43829;
	#10 counter$count = 43830;
	#10 counter$count = 43831;
	#10 counter$count = 43832;
	#10 counter$count = 43833;
	#10 counter$count = 43834;
	#10 counter$count = 43835;
	#10 counter$count = 43836;
	#10 counter$count = 43837;
	#10 counter$count = 43838;
	#10 counter$count = 43839;
	#10 counter$count = 43840;
	#10 counter$count = 43841;
	#10 counter$count = 43842;
	#10 counter$count = 43843;
	#10 counter$count = 43844;
	#10 counter$count = 43845;
	#10 counter$count = 43846;
	#10 counter$count = 43847;
	#10 counter$count = 43848;
	#10 counter$count = 43849;
	#10 counter$count = 43850;
	#10 counter$count = 43851;
	#10 counter$count = 43852;
	#10 counter$count = 43853;
	#10 counter$count = 43854;
	#10 counter$count = 43855;
	#10 counter$count = 43856;
	#10 counter$count = 43857;
	#10 counter$count = 43858;
	#10 counter$count = 43859;
	#10 counter$count = 43860;
	#10 counter$count = 43861;
	#10 counter$count = 43862;
	#10 counter$count = 43863;
	#10 counter$count = 43864;
	#10 counter$count = 43865;
	#10 counter$count = 43866;
	#10 counter$count = 43867;
	#10 counter$count = 43868;
	#10 counter$count = 43869;
	#10 counter$count = 43870;
	#10 counter$count = 43871;
	#10 counter$count = 43872;
	#10 counter$count = 43873;
	#10 counter$count = 43874;
	#10 counter$count = 43875;
	#10 counter$count = 43876;
	#10 counter$count = 43877;
	#10 counter$count = 43878;
	#10 counter$count = 43879;
	#10 counter$count = 43880;
	#10 counter$count = 43881;
	#10 counter$count = 43882;
	#10 counter$count = 43883;
	#10 counter$count = 43884;
	#10 counter$count = 43885;
	#10 counter$count = 43886;
	#10 counter$count = 43887;
	#10 counter$count = 43888;
	#10 counter$count = 43889;
	#10 counter$count = 43890;
	#10 counter$count = 43891;
	#10 counter$count = 43892;
	#10 counter$count = 43893;
	#10 counter$count = 43894;
	#10 counter$count = 43895;
	#10 counter$count = 43896;
	#10 counter$count = 43897;
	#10 counter$count = 43898;
	#10 counter$count = 43899;
	#10 counter$count = 43900;
	#10 counter$count = 43901;
	#10 counter$count = 43902;
	#10 counter$count = 43903;
	#10 counter$count = 43904;
	#10 counter$count = 43905;
	#10 counter$count = 43906;
	#10 counter$count = 43907;
	#10 counter$count = 43908;
	#10 counter$count = 43909;
	#10 counter$count = 43910;
	#10 counter$count = 43911;
	#10 counter$count = 43912;
	#10 counter$count = 43913;
	#10 counter$count = 43914;
	#10 counter$count = 43915;
	#10 counter$count = 43916;
	#10 counter$count = 43917;
	#10 counter$count = 43918;
	#10 counter$count = 43919;
	#10 counter$count = 43920;
	#10 counter$count = 43921;
	#10 counter$count = 43922;
	#10 counter$count = 43923;
	#10 counter$count = 43924;
	#10 counter$count = 43925;
	#10 counter$count = 43926;
	#10 counter$count = 43927;
	#10 counter$count = 43928;
	#10 counter$count = 43929;
	#10 counter$count = 43930;
	#10 counter$count = 43931;
	#10 counter$count = 43932;
	#10 counter$count = 43933;
	#10 counter$count = 43934;
	#10 counter$count = 43935;
	#10 counter$count = 43936;
	#10 counter$count = 43937;
	#10 counter$count = 43938;
	#10 counter$count = 43939;
	#10 counter$count = 43940;
	#10 counter$count = 43941;
	#10 counter$count = 43942;
	#10 counter$count = 43943;
	#10 counter$count = 43944;
	#10 counter$count = 43945;
	#10 counter$count = 43946;
	#10 counter$count = 43947;
	#10 counter$count = 43948;
	#10 counter$count = 43949;
	#10 counter$count = 43950;
	#10 counter$count = 43951;
	#10 counter$count = 43952;
	#10 counter$count = 43953;
	#10 counter$count = 43954;
	#10 counter$count = 43955;
	#10 counter$count = 43956;
	#10 counter$count = 43957;
	#10 counter$count = 43958;
	#10 counter$count = 43959;
	#10 counter$count = 43960;
	#10 counter$count = 43961;
	#10 counter$count = 43962;
	#10 counter$count = 43963;
	#10 counter$count = 43964;
	#10 counter$count = 43965;
	#10 counter$count = 43966;
	#10 counter$count = 43967;
	#10 counter$count = 43968;
	#10 counter$count = 43969;
	#10 counter$count = 43970;
	#10 counter$count = 43971;
	#10 counter$count = 43972;
	#10 counter$count = 43973;
	#10 counter$count = 43974;
	#10 counter$count = 43975;
	#10 counter$count = 43976;
	#10 counter$count = 43977;
	#10 counter$count = 43978;
	#10 counter$count = 43979;
	#10 counter$count = 43980;
	#10 counter$count = 43981;
	#10 counter$count = 43982;
	#10 counter$count = 43983;
	#10 counter$count = 43984;
	#10 counter$count = 43985;
	#10 counter$count = 43986;
	#10 counter$count = 43987;
	#10 counter$count = 43988;
	#10 counter$count = 43989;
	#10 counter$count = 43990;
	#10 counter$count = 43991;
	#10 counter$count = 43992;
	#10 counter$count = 43993;
	#10 counter$count = 43994;
	#10 counter$count = 43995;
	#10 counter$count = 43996;
	#10 counter$count = 43997;
	#10 counter$count = 43998;
	#10 counter$count = 43999;
	#10 counter$count = 44000;
	#10 counter$count = 44001;
	#10 counter$count = 44002;
	#10 counter$count = 44003;
	#10 counter$count = 44004;
	#10 counter$count = 44005;
	#10 counter$count = 44006;
	#10 counter$count = 44007;
	#10 counter$count = 44008;
	#10 counter$count = 44009;
	#10 counter$count = 44010;
	#10 counter$count = 44011;
	#10 counter$count = 44012;
	#10 counter$count = 44013;
	#10 counter$count = 44014;
	#10 counter$count = 44015;
	#10 counter$count = 44016;
	#10 counter$count = 44017;
	#10 counter$count = 44018;
	#10 counter$count = 44019;
	#10 counter$count = 44020;
	#10 counter$count = 44021;
	#10 counter$count = 44022;
	#10 counter$count = 44023;
	#10 counter$count = 44024;
	#10 counter$count = 44025;
	#10 counter$count = 44026;
	#10 counter$count = 44027;
	#10 counter$count = 44028;
	#10 counter$count = 44029;
	#10 counter$count = 44030;
	#10 counter$count = 44031;
	#10 counter$count = 44032;
	#10 counter$count = 44033;
	#10 counter$count = 44034;
	#10 counter$count = 44035;
	#10 counter$count = 44036;
	#10 counter$count = 44037;
	#10 counter$count = 44038;
	#10 counter$count = 44039;
	#10 counter$count = 44040;
	#10 counter$count = 44041;
	#10 counter$count = 44042;
	#10 counter$count = 44043;
	#10 counter$count = 44044;
	#10 counter$count = 44045;
	#10 counter$count = 44046;
	#10 counter$count = 44047;
	#10 counter$count = 44048;
	#10 counter$count = 44049;
	#10 counter$count = 44050;
	#10 counter$count = 44051;
	#10 counter$count = 44052;
	#10 counter$count = 44053;
	#10 counter$count = 44054;
	#10 counter$count = 44055;
	#10 counter$count = 44056;
	#10 counter$count = 44057;
	#10 counter$count = 44058;
	#10 counter$count = 44059;
	#10 counter$count = 44060;
	#10 counter$count = 44061;
	#10 counter$count = 44062;
	#10 counter$count = 44063;
	#10 counter$count = 44064;
	#10 counter$count = 44065;
	#10 counter$count = 44066;
	#10 counter$count = 44067;
	#10 counter$count = 44068;
	#10 counter$count = 44069;
	#10 counter$count = 44070;
	#10 counter$count = 44071;
	#10 counter$count = 44072;
	#10 counter$count = 44073;
	#10 counter$count = 44074;
	#10 counter$count = 44075;
	#10 counter$count = 44076;
	#10 counter$count = 44077;
	#10 counter$count = 44078;
	#10 counter$count = 44079;
	#10 counter$count = 44080;
	#10 counter$count = 44081;
	#10 counter$count = 44082;
	#10 counter$count = 44083;
	#10 counter$count = 44084;
	#10 counter$count = 44085;
	#10 counter$count = 44086;
	#10 counter$count = 44087;
	#10 counter$count = 44088;
	#10 counter$count = 44089;
	#10 counter$count = 44090;
	#10 counter$count = 44091;
	#10 counter$count = 44092;
	#10 counter$count = 44093;
	#10 counter$count = 44094;
	#10 counter$count = 44095;
	#10 counter$count = 44096;
	#10 counter$count = 44097;
	#10 counter$count = 44098;
	#10 counter$count = 44099;
	#10 counter$count = 44100;
	#10 counter$count = 44101;
	#10 counter$count = 44102;
	#10 counter$count = 44103;
	#10 counter$count = 44104;
	#10 counter$count = 44105;
	#10 counter$count = 44106;
	#10 counter$count = 44107;
	#10 counter$count = 44108;
	#10 counter$count = 44109;
	#10 counter$count = 44110;
	#10 counter$count = 44111;
	#10 counter$count = 44112;
	#10 counter$count = 44113;
	#10 counter$count = 44114;
	#10 counter$count = 44115;
	#10 counter$count = 44116;
	#10 counter$count = 44117;
	#10 counter$count = 44118;
	#10 counter$count = 44119;
	#10 counter$count = 44120;
	#10 counter$count = 44121;
	#10 counter$count = 44122;
	#10 counter$count = 44123;
	#10 counter$count = 44124;
	#10 counter$count = 44125;
	#10 counter$count = 44126;
	#10 counter$count = 44127;
	#10 counter$count = 44128;
	#10 counter$count = 44129;
	#10 counter$count = 44130;
	#10 counter$count = 44131;
	#10 counter$count = 44132;
	#10 counter$count = 44133;
	#10 counter$count = 44134;
	#10 counter$count = 44135;
	#10 counter$count = 44136;
	#10 counter$count = 44137;
	#10 counter$count = 44138;
	#10 counter$count = 44139;
	#10 counter$count = 44140;
	#10 counter$count = 44141;
	#10 counter$count = 44142;
	#10 counter$count = 44143;
	#10 counter$count = 44144;
	#10 counter$count = 44145;
	#10 counter$count = 44146;
	#10 counter$count = 44147;
	#10 counter$count = 44148;
	#10 counter$count = 44149;
	#10 counter$count = 44150;
	#10 counter$count = 44151;
	#10 counter$count = 44152;
	#10 counter$count = 44153;
	#10 counter$count = 44154;
	#10 counter$count = 44155;
	#10 counter$count = 44156;
	#10 counter$count = 44157;
	#10 counter$count = 44158;
	#10 counter$count = 44159;
	#10 counter$count = 44160;
	#10 counter$count = 44161;
	#10 counter$count = 44162;
	#10 counter$count = 44163;
	#10 counter$count = 44164;
	#10 counter$count = 44165;
	#10 counter$count = 44166;
	#10 counter$count = 44167;
	#10 counter$count = 44168;
	#10 counter$count = 44169;
	#10 counter$count = 44170;
	#10 counter$count = 44171;
	#10 counter$count = 44172;
	#10 counter$count = 44173;
	#10 counter$count = 44174;
	#10 counter$count = 44175;
	#10 counter$count = 44176;
	#10 counter$count = 44177;
	#10 counter$count = 44178;
	#10 counter$count = 44179;
	#10 counter$count = 44180;
	#10 counter$count = 44181;
	#10 counter$count = 44182;
	#10 counter$count = 44183;
	#10 counter$count = 44184;
	#10 counter$count = 44185;
	#10 counter$count = 44186;
	#10 counter$count = 44187;
	#10 counter$count = 44188;
	#10 counter$count = 44189;
	#10 counter$count = 44190;
	#10 counter$count = 44191;
	#10 counter$count = 44192;
	#10 counter$count = 44193;
	#10 counter$count = 44194;
	#10 counter$count = 44195;
	#10 counter$count = 44196;
	#10 counter$count = 44197;
	#10 counter$count = 44198;
	#10 counter$count = 44199;
	#10 counter$count = 44200;
	#10 counter$count = 44201;
	#10 counter$count = 44202;
	#10 counter$count = 44203;
	#10 counter$count = 44204;
	#10 counter$count = 44205;
	#10 counter$count = 44206;
	#10 counter$count = 44207;
	#10 counter$count = 44208;
	#10 counter$count = 44209;
	#10 counter$count = 44210;
	#10 counter$count = 44211;
	#10 counter$count = 44212;
	#10 counter$count = 44213;
	#10 counter$count = 44214;
	#10 counter$count = 44215;
	#10 counter$count = 44216;
	#10 counter$count = 44217;
	#10 counter$count = 44218;
	#10 counter$count = 44219;
	#10 counter$count = 44220;
	#10 counter$count = 44221;
	#10 counter$count = 44222;
	#10 counter$count = 44223;
	#10 counter$count = 44224;
	#10 counter$count = 44225;
	#10 counter$count = 44226;
	#10 counter$count = 44227;
	#10 counter$count = 44228;
	#10 counter$count = 44229;
	#10 counter$count = 44230;
	#10 counter$count = 44231;
	#10 counter$count = 44232;
	#10 counter$count = 44233;
	#10 counter$count = 44234;
	#10 counter$count = 44235;
	#10 counter$count = 44236;
	#10 counter$count = 44237;
	#10 counter$count = 44238;
	#10 counter$count = 44239;
	#10 counter$count = 44240;
	#10 counter$count = 44241;
	#10 counter$count = 44242;
	#10 counter$count = 44243;
	#10 counter$count = 44244;
	#10 counter$count = 44245;
	#10 counter$count = 44246;
	#10 counter$count = 44247;
	#10 counter$count = 44248;
	#10 counter$count = 44249;
	#10 counter$count = 44250;
	#10 counter$count = 44251;
	#10 counter$count = 44252;
	#10 counter$count = 44253;
	#10 counter$count = 44254;
	#10 counter$count = 44255;
	#10 counter$count = 44256;
	#10 counter$count = 44257;
	#10 counter$count = 44258;
	#10 counter$count = 44259;
	#10 counter$count = 44260;
	#10 counter$count = 44261;
	#10 counter$count = 44262;
	#10 counter$count = 44263;
	#10 counter$count = 44264;
	#10 counter$count = 44265;
	#10 counter$count = 44266;
	#10 counter$count = 44267;
	#10 counter$count = 44268;
	#10 counter$count = 44269;
	#10 counter$count = 44270;
	#10 counter$count = 44271;
	#10 counter$count = 44272;
	#10 counter$count = 44273;
	#10 counter$count = 44274;
	#10 counter$count = 44275;
	#10 counter$count = 44276;
	#10 counter$count = 44277;
	#10 counter$count = 44278;
	#10 counter$count = 44279;
	#10 counter$count = 44280;
	#10 counter$count = 44281;
	#10 counter$count = 44282;
	#10 counter$count = 44283;
	#10 counter$count = 44284;
	#10 counter$count = 44285;
	#10 counter$count = 44286;
	#10 counter$count = 44287;
	#10 counter$count = 44288;
	#10 counter$count = 44289;
	#10 counter$count = 44290;
	#10 counter$count = 44291;
	#10 counter$count = 44292;
	#10 counter$count = 44293;
	#10 counter$count = 44294;
	#10 counter$count = 44295;
	#10 counter$count = 44296;
	#10 counter$count = 44297;
	#10 counter$count = 44298;
	#10 counter$count = 44299;
	#10 counter$count = 44300;
	#10 counter$count = 44301;
	#10 counter$count = 44302;
	#10 counter$count = 44303;
	#10 counter$count = 44304;
	#10 counter$count = 44305;
	#10 counter$count = 44306;
	#10 counter$count = 44307;
	#10 counter$count = 44308;
	#10 counter$count = 44309;
	#10 counter$count = 44310;
	#10 counter$count = 44311;
	#10 counter$count = 44312;
	#10 counter$count = 44313;
	#10 counter$count = 44314;
	#10 counter$count = 44315;
	#10 counter$count = 44316;
	#10 counter$count = 44317;
	#10 counter$count = 44318;
	#10 counter$count = 44319;
	#10 counter$count = 44320;
	#10 counter$count = 44321;
	#10 counter$count = 44322;
	#10 counter$count = 44323;
	#10 counter$count = 44324;
	#10 counter$count = 44325;
	#10 counter$count = 44326;
	#10 counter$count = 44327;
	#10 counter$count = 44328;
	#10 counter$count = 44329;
	#10 counter$count = 44330;
	#10 counter$count = 44331;
	#10 counter$count = 44332;
	#10 counter$count = 44333;
	#10 counter$count = 44334;
	#10 counter$count = 44335;
	#10 counter$count = 44336;
	#10 counter$count = 44337;
	#10 counter$count = 44338;
	#10 counter$count = 44339;
	#10 counter$count = 44340;
	#10 counter$count = 44341;
	#10 counter$count = 44342;
	#10 counter$count = 44343;
	#10 counter$count = 44344;
	#10 counter$count = 44345;
	#10 counter$count = 44346;
	#10 counter$count = 44347;
	#10 counter$count = 44348;
	#10 counter$count = 44349;
	#10 counter$count = 44350;
	#10 counter$count = 44351;
	#10 counter$count = 44352;
	#10 counter$count = 44353;
	#10 counter$count = 44354;
	#10 counter$count = 44355;
	#10 counter$count = 44356;
	#10 counter$count = 44357;
	#10 counter$count = 44358;
	#10 counter$count = 44359;
	#10 counter$count = 44360;
	#10 counter$count = 44361;
	#10 counter$count = 44362;
	#10 counter$count = 44363;
	#10 counter$count = 44364;
	#10 counter$count = 44365;
	#10 counter$count = 44366;
	#10 counter$count = 44367;
	#10 counter$count = 44368;
	#10 counter$count = 44369;
	#10 counter$count = 44370;
	#10 counter$count = 44371;
	#10 counter$count = 44372;
	#10 counter$count = 44373;
	#10 counter$count = 44374;
	#10 counter$count = 44375;
	#10 counter$count = 44376;
	#10 counter$count = 44377;
	#10 counter$count = 44378;
	#10 counter$count = 44379;
	#10 counter$count = 44380;
	#10 counter$count = 44381;
	#10 counter$count = 44382;
	#10 counter$count = 44383;
	#10 counter$count = 44384;
	#10 counter$count = 44385;
	#10 counter$count = 44386;
	#10 counter$count = 44387;
	#10 counter$count = 44388;
	#10 counter$count = 44389;
	#10 counter$count = 44390;
	#10 counter$count = 44391;
	#10 counter$count = 44392;
	#10 counter$count = 44393;
	#10 counter$count = 44394;
	#10 counter$count = 44395;
	#10 counter$count = 44396;
	#10 counter$count = 44397;
	#10 counter$count = 44398;
	#10 counter$count = 44399;
	#10 counter$count = 44400;
	#10 counter$count = 44401;
	#10 counter$count = 44402;
	#10 counter$count = 44403;
	#10 counter$count = 44404;
	#10 counter$count = 44405;
	#10 counter$count = 44406;
	#10 counter$count = 44407;
	#10 counter$count = 44408;
	#10 counter$count = 44409;
	#10 counter$count = 44410;
	#10 counter$count = 44411;
	#10 counter$count = 44412;
	#10 counter$count = 44413;
	#10 counter$count = 44414;
	#10 counter$count = 44415;
	#10 counter$count = 44416;
	#10 counter$count = 44417;
	#10 counter$count = 44418;
	#10 counter$count = 44419;
	#10 counter$count = 44420;
	#10 counter$count = 44421;
	#10 counter$count = 44422;
	#10 counter$count = 44423;
	#10 counter$count = 44424;
	#10 counter$count = 44425;
	#10 counter$count = 44426;
	#10 counter$count = 44427;
	#10 counter$count = 44428;
	#10 counter$count = 44429;
	#10 counter$count = 44430;
	#10 counter$count = 44431;
	#10 counter$count = 44432;
	#10 counter$count = 44433;
	#10 counter$count = 44434;
	#10 counter$count = 44435;
	#10 counter$count = 44436;
	#10 counter$count = 44437;
	#10 counter$count = 44438;
	#10 counter$count = 44439;
	#10 counter$count = 44440;
	#10 counter$count = 44441;
	#10 counter$count = 44442;
	#10 counter$count = 44443;
	#10 counter$count = 44444;
	#10 counter$count = 44445;
	#10 counter$count = 44446;
	#10 counter$count = 44447;
	#10 counter$count = 44448;
	#10 counter$count = 44449;
	#10 counter$count = 44450;
	#10 counter$count = 44451;
	#10 counter$count = 44452;
	#10 counter$count = 44453;
	#10 counter$count = 44454;
	#10 counter$count = 44455;
	#10 counter$count = 44456;
	#10 counter$count = 44457;
	#10 counter$count = 44458;
	#10 counter$count = 44459;
	#10 counter$count = 44460;
	#10 counter$count = 44461;
	#10 counter$count = 44462;
	#10 counter$count = 44463;
	#10 counter$count = 44464;
	#10 counter$count = 44465;
	#10 counter$count = 44466;
	#10 counter$count = 44467;
	#10 counter$count = 44468;
	#10 counter$count = 44469;
	#10 counter$count = 44470;
	#10 counter$count = 44471;
	#10 counter$count = 44472;
	#10 counter$count = 44473;
	#10 counter$count = 44474;
	#10 counter$count = 44475;
	#10 counter$count = 44476;
	#10 counter$count = 44477;
	#10 counter$count = 44478;
	#10 counter$count = 44479;
	#10 counter$count = 44480;
	#10 counter$count = 44481;
	#10 counter$count = 44482;
	#10 counter$count = 44483;
	#10 counter$count = 44484;
	#10 counter$count = 44485;
	#10 counter$count = 44486;
	#10 counter$count = 44487;
	#10 counter$count = 44488;
	#10 counter$count = 44489;
	#10 counter$count = 44490;
	#10 counter$count = 44491;
	#10 counter$count = 44492;
	#10 counter$count = 44493;
	#10 counter$count = 44494;
	#10 counter$count = 44495;
	#10 counter$count = 44496;
	#10 counter$count = 44497;
	#10 counter$count = 44498;
	#10 counter$count = 44499;
	#10 counter$count = 44500;
	#10 counter$count = 44501;
	#10 counter$count = 44502;
	#10 counter$count = 44503;
	#10 counter$count = 44504;
	#10 counter$count = 44505;
	#10 counter$count = 44506;
	#10 counter$count = 44507;
	#10 counter$count = 44508;
	#10 counter$count = 44509;
	#10 counter$count = 44510;
	#10 counter$count = 44511;
	#10 counter$count = 44512;
	#10 counter$count = 44513;
	#10 counter$count = 44514;
	#10 counter$count = 44515;
	#10 counter$count = 44516;
	#10 counter$count = 44517;
	#10 counter$count = 44518;
	#10 counter$count = 44519;
	#10 counter$count = 44520;
	#10 counter$count = 44521;
	#10 counter$count = 44522;
	#10 counter$count = 44523;
	#10 counter$count = 44524;
	#10 counter$count = 44525;
	#10 counter$count = 44526;
	#10 counter$count = 44527;
	#10 counter$count = 44528;
	#10 counter$count = 44529;
	#10 counter$count = 44530;
	#10 counter$count = 44531;
	#10 counter$count = 44532;
	#10 counter$count = 44533;
	#10 counter$count = 44534;
	#10 counter$count = 44535;
	#10 counter$count = 44536;
	#10 counter$count = 44537;
	#10 counter$count = 44538;
	#10 counter$count = 44539;
	#10 counter$count = 44540;
	#10 counter$count = 44541;
	#10 counter$count = 44542;
	#10 counter$count = 44543;
	#10 counter$count = 44544;
	#10 counter$count = 44545;
	#10 counter$count = 44546;
	#10 counter$count = 44547;
	#10 counter$count = 44548;
	#10 counter$count = 44549;
	#10 counter$count = 44550;
	#10 counter$count = 44551;
	#10 counter$count = 44552;
	#10 counter$count = 44553;
	#10 counter$count = 44554;
	#10 counter$count = 44555;
	#10 counter$count = 44556;
	#10 counter$count = 44557;
	#10 counter$count = 44558;
	#10 counter$count = 44559;
	#10 counter$count = 44560;
	#10 counter$count = 44561;
	#10 counter$count = 44562;
	#10 counter$count = 44563;
	#10 counter$count = 44564;
	#10 counter$count = 44565;
	#10 counter$count = 44566;
	#10 counter$count = 44567;
	#10 counter$count = 44568;
	#10 counter$count = 44569;
	#10 counter$count = 44570;
	#10 counter$count = 44571;
	#10 counter$count = 44572;
	#10 counter$count = 44573;
	#10 counter$count = 44574;
	#10 counter$count = 44575;
	#10 counter$count = 44576;
	#10 counter$count = 44577;
	#10 counter$count = 44578;
	#10 counter$count = 44579;
	#10 counter$count = 44580;
	#10 counter$count = 44581;
	#10 counter$count = 44582;
	#10 counter$count = 44583;
	#10 counter$count = 44584;
	#10 counter$count = 44585;
	#10 counter$count = 44586;
	#10 counter$count = 44587;
	#10 counter$count = 44588;
	#10 counter$count = 44589;
	#10 counter$count = 44590;
	#10 counter$count = 44591;
	#10 counter$count = 44592;
	#10 counter$count = 44593;
	#10 counter$count = 44594;
	#10 counter$count = 44595;
	#10 counter$count = 44596;
	#10 counter$count = 44597;
	#10 counter$count = 44598;
	#10 counter$count = 44599;
	#10 counter$count = 44600;
	#10 counter$count = 44601;
	#10 counter$count = 44602;
	#10 counter$count = 44603;
	#10 counter$count = 44604;
	#10 counter$count = 44605;
	#10 counter$count = 44606;
	#10 counter$count = 44607;
	#10 counter$count = 44608;
	#10 counter$count = 44609;
	#10 counter$count = 44610;
	#10 counter$count = 44611;
	#10 counter$count = 44612;
	#10 counter$count = 44613;
	#10 counter$count = 44614;
	#10 counter$count = 44615;
	#10 counter$count = 44616;
	#10 counter$count = 44617;
	#10 counter$count = 44618;
	#10 counter$count = 44619;
	#10 counter$count = 44620;
	#10 counter$count = 44621;
	#10 counter$count = 44622;
	#10 counter$count = 44623;
	#10 counter$count = 44624;
	#10 counter$count = 44625;
	#10 counter$count = 44626;
	#10 counter$count = 44627;
	#10 counter$count = 44628;
	#10 counter$count = 44629;
	#10 counter$count = 44630;
	#10 counter$count = 44631;
	#10 counter$count = 44632;
	#10 counter$count = 44633;
	#10 counter$count = 44634;
	#10 counter$count = 44635;
	#10 counter$count = 44636;
	#10 counter$count = 44637;
	#10 counter$count = 44638;
	#10 counter$count = 44639;
	#10 counter$count = 44640;
	#10 counter$count = 44641;
	#10 counter$count = 44642;
	#10 counter$count = 44643;
	#10 counter$count = 44644;
	#10 counter$count = 44645;
	#10 counter$count = 44646;
	#10 counter$count = 44647;
	#10 counter$count = 44648;
	#10 counter$count = 44649;
	#10 counter$count = 44650;
	#10 counter$count = 44651;
	#10 counter$count = 44652;
	#10 counter$count = 44653;
	#10 counter$count = 44654;
	#10 counter$count = 44655;
	#10 counter$count = 44656;
	#10 counter$count = 44657;
	#10 counter$count = 44658;
	#10 counter$count = 44659;
	#10 counter$count = 44660;
	#10 counter$count = 44661;
	#10 counter$count = 44662;
	#10 counter$count = 44663;
	#10 counter$count = 44664;
	#10 counter$count = 44665;
	#10 counter$count = 44666;
	#10 counter$count = 44667;
	#10 counter$count = 44668;
	#10 counter$count = 44669;
	#10 counter$count = 44670;
	#10 counter$count = 44671;
	#10 counter$count = 44672;
	#10 counter$count = 44673;
	#10 counter$count = 44674;
	#10 counter$count = 44675;
	#10 counter$count = 44676;
	#10 counter$count = 44677;
	#10 counter$count = 44678;
	#10 counter$count = 44679;
	#10 counter$count = 44680;
	#10 counter$count = 44681;
	#10 counter$count = 44682;
	#10 counter$count = 44683;
	#10 counter$count = 44684;
	#10 counter$count = 44685;
	#10 counter$count = 44686;
	#10 counter$count = 44687;
	#10 counter$count = 44688;
	#10 counter$count = 44689;
	#10 counter$count = 44690;
	#10 counter$count = 44691;
	#10 counter$count = 44692;
	#10 counter$count = 44693;
	#10 counter$count = 44694;
	#10 counter$count = 44695;
	#10 counter$count = 44696;
	#10 counter$count = 44697;
	#10 counter$count = 44698;
	#10 counter$count = 44699;
	#10 counter$count = 44700;
	#10 counter$count = 44701;
	#10 counter$count = 44702;
	#10 counter$count = 44703;
	#10 counter$count = 44704;
	#10 counter$count = 44705;
	#10 counter$count = 44706;
	#10 counter$count = 44707;
	#10 counter$count = 44708;
	#10 counter$count = 44709;
	#10 counter$count = 44710;
	#10 counter$count = 44711;
	#10 counter$count = 44712;
	#10 counter$count = 44713;
	#10 counter$count = 44714;
	#10 counter$count = 44715;
	#10 counter$count = 44716;
	#10 counter$count = 44717;
	#10 counter$count = 44718;
	#10 counter$count = 44719;
	#10 counter$count = 44720;
	#10 counter$count = 44721;
	#10 counter$count = 44722;
	#10 counter$count = 44723;
	#10 counter$count = 44724;
	#10 counter$count = 44725;
	#10 counter$count = 44726;
	#10 counter$count = 44727;
	#10 counter$count = 44728;
	#10 counter$count = 44729;
	#10 counter$count = 44730;
	#10 counter$count = 44731;
	#10 counter$count = 44732;
	#10 counter$count = 44733;
	#10 counter$count = 44734;
	#10 counter$count = 44735;
	#10 counter$count = 44736;
	#10 counter$count = 44737;
	#10 counter$count = 44738;
	#10 counter$count = 44739;
	#10 counter$count = 44740;
	#10 counter$count = 44741;
	#10 counter$count = 44742;
	#10 counter$count = 44743;
	#10 counter$count = 44744;
	#10 counter$count = 44745;
	#10 counter$count = 44746;
	#10 counter$count = 44747;
	#10 counter$count = 44748;
	#10 counter$count = 44749;
	#10 counter$count = 44750;
	#10 counter$count = 44751;
	#10 counter$count = 44752;
	#10 counter$count = 44753;
	#10 counter$count = 44754;
	#10 counter$count = 44755;
	#10 counter$count = 44756;
	#10 counter$count = 44757;
	#10 counter$count = 44758;
	#10 counter$count = 44759;
	#10 counter$count = 44760;
	#10 counter$count = 44761;
	#10 counter$count = 44762;
	#10 counter$count = 44763;
	#10 counter$count = 44764;
	#10 counter$count = 44765;
	#10 counter$count = 44766;
	#10 counter$count = 44767;
	#10 counter$count = 44768;
	#10 counter$count = 44769;
	#10 counter$count = 44770;
	#10 counter$count = 44771;
	#10 counter$count = 44772;
	#10 counter$count = 44773;
	#10 counter$count = 44774;
	#10 counter$count = 44775;
	#10 counter$count = 44776;
	#10 counter$count = 44777;
	#10 counter$count = 44778;
	#10 counter$count = 44779;
	#10 counter$count = 44780;
	#10 counter$count = 44781;
	#10 counter$count = 44782;
	#10 counter$count = 44783;
	#10 counter$count = 44784;
	#10 counter$count = 44785;
	#10 counter$count = 44786;
	#10 counter$count = 44787;
	#10 counter$count = 44788;
	#10 counter$count = 44789;
	#10 counter$count = 44790;
	#10 counter$count = 44791;
	#10 counter$count = 44792;
	#10 counter$count = 44793;
	#10 counter$count = 44794;
	#10 counter$count = 44795;
	#10 counter$count = 44796;
	#10 counter$count = 44797;
	#10 counter$count = 44798;
	#10 counter$count = 44799;
	#10 counter$count = 44800;
	#10 counter$count = 44801;
	#10 counter$count = 44802;
	#10 counter$count = 44803;
	#10 counter$count = 44804;
	#10 counter$count = 44805;
	#10 counter$count = 44806;
	#10 counter$count = 44807;
	#10 counter$count = 44808;
	#10 counter$count = 44809;
	#10 counter$count = 44810;
	#10 counter$count = 44811;
	#10 counter$count = 44812;
	#10 counter$count = 44813;
	#10 counter$count = 44814;
	#10 counter$count = 44815;
	#10 counter$count = 44816;
	#10 counter$count = 44817;
	#10 counter$count = 44818;
	#10 counter$count = 44819;
	#10 counter$count = 44820;
	#10 counter$count = 44821;
	#10 counter$count = 44822;
	#10 counter$count = 44823;
	#10 counter$count = 44824;
	#10 counter$count = 44825;
	#10 counter$count = 44826;
	#10 counter$count = 44827;
	#10 counter$count = 44828;
	#10 counter$count = 44829;
	#10 counter$count = 44830;
	#10 counter$count = 44831;
	#10 counter$count = 44832;
	#10 counter$count = 44833;
	#10 counter$count = 44834;
	#10 counter$count = 44835;
	#10 counter$count = 44836;
	#10 counter$count = 44837;
	#10 counter$count = 44838;
	#10 counter$count = 44839;
	#10 counter$count = 44840;
	#10 counter$count = 44841;
	#10 counter$count = 44842;
	#10 counter$count = 44843;
	#10 counter$count = 44844;
	#10 counter$count = 44845;
	#10 counter$count = 44846;
	#10 counter$count = 44847;
	#10 counter$count = 44848;
	#10 counter$count = 44849;
	#10 counter$count = 44850;
	#10 counter$count = 44851;
	#10 counter$count = 44852;
	#10 counter$count = 44853;
	#10 counter$count = 44854;
	#10 counter$count = 44855;
	#10 counter$count = 44856;
	#10 counter$count = 44857;
	#10 counter$count = 44858;
	#10 counter$count = 44859;
	#10 counter$count = 44860;
	#10 counter$count = 44861;
	#10 counter$count = 44862;
	#10 counter$count = 44863;
	#10 counter$count = 44864;
	#10 counter$count = 44865;
	#10 counter$count = 44866;
	#10 counter$count = 44867;
	#10 counter$count = 44868;
	#10 counter$count = 44869;
	#10 counter$count = 44870;
	#10 counter$count = 44871;
	#10 counter$count = 44872;
	#10 counter$count = 44873;
	#10 counter$count = 44874;
	#10 counter$count = 44875;
	#10 counter$count = 44876;
	#10 counter$count = 44877;
	#10 counter$count = 44878;
	#10 counter$count = 44879;
	#10 counter$count = 44880;
	#10 counter$count = 44881;
	#10 counter$count = 44882;
	#10 counter$count = 44883;
	#10 counter$count = 44884;
	#10 counter$count = 44885;
	#10 counter$count = 44886;
	#10 counter$count = 44887;
	#10 counter$count = 44888;
	#10 counter$count = 44889;
	#10 counter$count = 44890;
	#10 counter$count = 44891;
	#10 counter$count = 44892;
	#10 counter$count = 44893;
	#10 counter$count = 44894;
	#10 counter$count = 44895;
	#10 counter$count = 44896;
	#10 counter$count = 44897;
	#10 counter$count = 44898;
	#10 counter$count = 44899;
	#10 counter$count = 44900;
	#10 counter$count = 44901;
	#10 counter$count = 44902;
	#10 counter$count = 44903;
	#10 counter$count = 44904;
	#10 counter$count = 44905;
	#10 counter$count = 44906;
	#10 counter$count = 44907;
	#10 counter$count = 44908;
	#10 counter$count = 44909;
	#10 counter$count = 44910;
	#10 counter$count = 44911;
	#10 counter$count = 44912;
	#10 counter$count = 44913;
	#10 counter$count = 44914;
	#10 counter$count = 44915;
	#10 counter$count = 44916;
	#10 counter$count = 44917;
	#10 counter$count = 44918;
	#10 counter$count = 44919;
	#10 counter$count = 44920;
	#10 counter$count = 44921;
	#10 counter$count = 44922;
	#10 counter$count = 44923;
	#10 counter$count = 44924;
	#10 counter$count = 44925;
	#10 counter$count = 44926;
	#10 counter$count = 44927;
	#10 counter$count = 44928;
	#10 counter$count = 44929;
	#10 counter$count = 44930;
	#10 counter$count = 44931;
	#10 counter$count = 44932;
	#10 counter$count = 44933;
	#10 counter$count = 44934;
	#10 counter$count = 44935;
	#10 counter$count = 44936;
	#10 counter$count = 44937;
	#10 counter$count = 44938;
	#10 counter$count = 44939;
	#10 counter$count = 44940;
	#10 counter$count = 44941;
	#10 counter$count = 44942;
	#10 counter$count = 44943;
	#10 counter$count = 44944;
	#10 counter$count = 44945;
	#10 counter$count = 44946;
	#10 counter$count = 44947;
	#10 counter$count = 44948;
	#10 counter$count = 44949;
	#10 counter$count = 44950;
	#10 counter$count = 44951;
	#10 counter$count = 44952;
	#10 counter$count = 44953;
	#10 counter$count = 44954;
	#10 counter$count = 44955;
	#10 counter$count = 44956;
	#10 counter$count = 44957;
	#10 counter$count = 44958;
	#10 counter$count = 44959;
	#10 counter$count = 44960;
	#10 counter$count = 44961;
	#10 counter$count = 44962;
	#10 counter$count = 44963;
	#10 counter$count = 44964;
	#10 counter$count = 44965;
	#10 counter$count = 44966;
	#10 counter$count = 44967;
	#10 counter$count = 44968;
	#10 counter$count = 44969;
	#10 counter$count = 44970;
	#10 counter$count = 44971;
	#10 counter$count = 44972;
	#10 counter$count = 44973;
	#10 counter$count = 44974;
	#10 counter$count = 44975;
	#10 counter$count = 44976;
	#10 counter$count = 44977;
	#10 counter$count = 44978;
	#10 counter$count = 44979;
	#10 counter$count = 44980;
	#10 counter$count = 44981;
	#10 counter$count = 44982;
	#10 counter$count = 44983;
	#10 counter$count = 44984;
	#10 counter$count = 44985;
	#10 counter$count = 44986;
	#10 counter$count = 44987;
	#10 counter$count = 44988;
	#10 counter$count = 44989;
	#10 counter$count = 44990;
	#10 counter$count = 44991;
	#10 counter$count = 44992;
	#10 counter$count = 44993;
	#10 counter$count = 44994;
	#10 counter$count = 44995;
	#10 counter$count = 44996;
	#10 counter$count = 44997;
	#10 counter$count = 44998;
	#10 counter$count = 44999;
	#10 counter$count = 45000;
	#10 counter$count = 45001;
	#10 counter$count = 45002;
	#10 counter$count = 45003;
	#10 counter$count = 45004;
	#10 counter$count = 45005;
	#10 counter$count = 45006;
	#10 counter$count = 45007;
	#10 counter$count = 45008;
	#10 counter$count = 45009;
	#10 counter$count = 45010;
	#10 counter$count = 45011;
	#10 counter$count = 45012;
	#10 counter$count = 45013;
	#10 counter$count = 45014;
	#10 counter$count = 45015;
	#10 counter$count = 45016;
	#10 counter$count = 45017;
	#10 counter$count = 45018;
	#10 counter$count = 45019;
	#10 counter$count = 45020;
	#10 counter$count = 45021;
	#10 counter$count = 45022;
	#10 counter$count = 45023;
	#10 counter$count = 45024;
	#10 counter$count = 45025;
	#10 counter$count = 45026;
	#10 counter$count = 45027;
	#10 counter$count = 45028;
	#10 counter$count = 45029;
	#10 counter$count = 45030;
	#10 counter$count = 45031;
	#10 counter$count = 45032;
	#10 counter$count = 45033;
	#10 counter$count = 45034;
	#10 counter$count = 45035;
	#10 counter$count = 45036;
	#10 counter$count = 45037;
	#10 counter$count = 45038;
	#10 counter$count = 45039;
	#10 counter$count = 45040;
	#10 counter$count = 45041;
	#10 counter$count = 45042;
	#10 counter$count = 45043;
	#10 counter$count = 45044;
	#10 counter$count = 45045;
	#10 counter$count = 45046;
	#10 counter$count = 45047;
	#10 counter$count = 45048;
	#10 counter$count = 45049;
	#10 counter$count = 45050;
	#10 counter$count = 45051;
	#10 counter$count = 45052;
	#10 counter$count = 45053;
	#10 counter$count = 45054;
	#10 counter$count = 45055;
	#10 counter$count = 45056;
	#10 counter$count = 45057;
	#10 counter$count = 45058;
	#10 counter$count = 45059;
	#10 counter$count = 45060;
	#10 counter$count = 45061;
	#10 counter$count = 45062;
	#10 counter$count = 45063;
	#10 counter$count = 45064;
	#10 counter$count = 45065;
	#10 counter$count = 45066;
	#10 counter$count = 45067;
	#10 counter$count = 45068;
	#10 counter$count = 45069;
	#10 counter$count = 45070;
	#10 counter$count = 45071;
	#10 counter$count = 45072;
	#10 counter$count = 45073;
	#10 counter$count = 45074;
	#10 counter$count = 45075;
	#10 counter$count = 45076;
	#10 counter$count = 45077;
	#10 counter$count = 45078;
	#10 counter$count = 45079;
	#10 counter$count = 45080;
	#10 counter$count = 45081;
	#10 counter$count = 45082;
	#10 counter$count = 45083;
	#10 counter$count = 45084;
	#10 counter$count = 45085;
	#10 counter$count = 45086;
	#10 counter$count = 45087;
	#10 counter$count = 45088;
	#10 counter$count = 45089;
	#10 counter$count = 45090;
	#10 counter$count = 45091;
	#10 counter$count = 45092;
	#10 counter$count = 45093;
	#10 counter$count = 45094;
	#10 counter$count = 45095;
	#10 counter$count = 45096;
	#10 counter$count = 45097;
	#10 counter$count = 45098;
	#10 counter$count = 45099;
	#10 counter$count = 45100;
	#10 counter$count = 45101;
	#10 counter$count = 45102;
	#10 counter$count = 45103;
	#10 counter$count = 45104;
	#10 counter$count = 45105;
	#10 counter$count = 45106;
	#10 counter$count = 45107;
	#10 counter$count = 45108;
	#10 counter$count = 45109;
	#10 counter$count = 45110;
	#10 counter$count = 45111;
	#10 counter$count = 45112;
	#10 counter$count = 45113;
	#10 counter$count = 45114;
	#10 counter$count = 45115;
	#10 counter$count = 45116;
	#10 counter$count = 45117;
	#10 counter$count = 45118;
	#10 counter$count = 45119;
	#10 counter$count = 45120;
	#10 counter$count = 45121;
	#10 counter$count = 45122;
	#10 counter$count = 45123;
	#10 counter$count = 45124;
	#10 counter$count = 45125;
	#10 counter$count = 45126;
	#10 counter$count = 45127;
	#10 counter$count = 45128;
	#10 counter$count = 45129;
	#10 counter$count = 45130;
	#10 counter$count = 45131;
	#10 counter$count = 45132;
	#10 counter$count = 45133;
	#10 counter$count = 45134;
	#10 counter$count = 45135;
	#10 counter$count = 45136;
	#10 counter$count = 45137;
	#10 counter$count = 45138;
	#10 counter$count = 45139;
	#10 counter$count = 45140;
	#10 counter$count = 45141;
	#10 counter$count = 45142;
	#10 counter$count = 45143;
	#10 counter$count = 45144;
	#10 counter$count = 45145;
	#10 counter$count = 45146;
	#10 counter$count = 45147;
	#10 counter$count = 45148;
	#10 counter$count = 45149;
	#10 counter$count = 45150;
	#10 counter$count = 45151;
	#10 counter$count = 45152;
	#10 counter$count = 45153;
	#10 counter$count = 45154;
	#10 counter$count = 45155;
	#10 counter$count = 45156;
	#10 counter$count = 45157;
	#10 counter$count = 45158;
	#10 counter$count = 45159;
	#10 counter$count = 45160;
	#10 counter$count = 45161;
	#10 counter$count = 45162;
	#10 counter$count = 45163;
	#10 counter$count = 45164;
	#10 counter$count = 45165;
	#10 counter$count = 45166;
	#10 counter$count = 45167;
	#10 counter$count = 45168;
	#10 counter$count = 45169;
	#10 counter$count = 45170;
	#10 counter$count = 45171;
	#10 counter$count = 45172;
	#10 counter$count = 45173;
	#10 counter$count = 45174;
	#10 counter$count = 45175;
	#10 counter$count = 45176;
	#10 counter$count = 45177;
	#10 counter$count = 45178;
	#10 counter$count = 45179;
	#10 counter$count = 45180;
	#10 counter$count = 45181;
	#10 counter$count = 45182;
	#10 counter$count = 45183;
	#10 counter$count = 45184;
	#10 counter$count = 45185;
	#10 counter$count = 45186;
	#10 counter$count = 45187;
	#10 counter$count = 45188;
	#10 counter$count = 45189;
	#10 counter$count = 45190;
	#10 counter$count = 45191;
	#10 counter$count = 45192;
	#10 counter$count = 45193;
	#10 counter$count = 45194;
	#10 counter$count = 45195;
	#10 counter$count = 45196;
	#10 counter$count = 45197;
	#10 counter$count = 45198;
	#10 counter$count = 45199;
	#10 counter$count = 45200;
	#10 counter$count = 45201;
	#10 counter$count = 45202;
	#10 counter$count = 45203;
	#10 counter$count = 45204;
	#10 counter$count = 45205;
	#10 counter$count = 45206;
	#10 counter$count = 45207;
	#10 counter$count = 45208;
	#10 counter$count = 45209;
	#10 counter$count = 45210;
	#10 counter$count = 45211;
	#10 counter$count = 45212;
	#10 counter$count = 45213;
	#10 counter$count = 45214;
	#10 counter$count = 45215;
	#10 counter$count = 45216;
	#10 counter$count = 45217;
	#10 counter$count = 45218;
	#10 counter$count = 45219;
	#10 counter$count = 45220;
	#10 counter$count = 45221;
	#10 counter$count = 45222;
	#10 counter$count = 45223;
	#10 counter$count = 45224;
	#10 counter$count = 45225;
	#10 counter$count = 45226;
	#10 counter$count = 45227;
	#10 counter$count = 45228;
	#10 counter$count = 45229;
	#10 counter$count = 45230;
	#10 counter$count = 45231;
	#10 counter$count = 45232;
	#10 counter$count = 45233;
	#10 counter$count = 45234;
	#10 counter$count = 45235;
	#10 counter$count = 45236;
	#10 counter$count = 45237;
	#10 counter$count = 45238;
	#10 counter$count = 45239;
	#10 counter$count = 45240;
	#10 counter$count = 45241;
	#10 counter$count = 45242;
	#10 counter$count = 45243;
	#10 counter$count = 45244;
	#10 counter$count = 45245;
	#10 counter$count = 45246;
	#10 counter$count = 45247;
	#10 counter$count = 45248;
	#10 counter$count = 45249;
	#10 counter$count = 45250;
	#10 counter$count = 45251;
	#10 counter$count = 45252;
	#10 counter$count = 45253;
	#10 counter$count = 45254;
	#10 counter$count = 45255;
	#10 counter$count = 45256;
	#10 counter$count = 45257;
	#10 counter$count = 45258;
	#10 counter$count = 45259;
	#10 counter$count = 45260;
	#10 counter$count = 45261;
	#10 counter$count = 45262;
	#10 counter$count = 45263;
	#10 counter$count = 45264;
	#10 counter$count = 45265;
	#10 counter$count = 45266;
	#10 counter$count = 45267;
	#10 counter$count = 45268;
	#10 counter$count = 45269;
	#10 counter$count = 45270;
	#10 counter$count = 45271;
	#10 counter$count = 45272;
	#10 counter$count = 45273;
	#10 counter$count = 45274;
	#10 counter$count = 45275;
	#10 counter$count = 45276;
	#10 counter$count = 45277;
	#10 counter$count = 45278;
	#10 counter$count = 45279;
	#10 counter$count = 45280;
	#10 counter$count = 45281;
	#10 counter$count = 45282;
	#10 counter$count = 45283;
	#10 counter$count = 45284;
	#10 counter$count = 45285;
	#10 counter$count = 45286;
	#10 counter$count = 45287;
	#10 counter$count = 45288;
	#10 counter$count = 45289;
	#10 counter$count = 45290;
	#10 counter$count = 45291;
	#10 counter$count = 45292;
	#10 counter$count = 45293;
	#10 counter$count = 45294;
	#10 counter$count = 45295;
	#10 counter$count = 45296;
	#10 counter$count = 45297;
	#10 counter$count = 45298;
	#10 counter$count = 45299;
	#10 counter$count = 45300;
	#10 counter$count = 45301;
	#10 counter$count = 45302;
	#10 counter$count = 45303;
	#10 counter$count = 45304;
	#10 counter$count = 45305;
	#10 counter$count = 45306;
	#10 counter$count = 45307;
	#10 counter$count = 45308;
	#10 counter$count = 45309;
	#10 counter$count = 45310;
	#10 counter$count = 45311;
	#10 counter$count = 45312;
	#10 counter$count = 45313;
	#10 counter$count = 45314;
	#10 counter$count = 45315;
	#10 counter$count = 45316;
	#10 counter$count = 45317;
	#10 counter$count = 45318;
	#10 counter$count = 45319;
	#10 counter$count = 45320;
	#10 counter$count = 45321;
	#10 counter$count = 45322;
	#10 counter$count = 45323;
	#10 counter$count = 45324;
	#10 counter$count = 45325;
	#10 counter$count = 45326;
	#10 counter$count = 45327;
	#10 counter$count = 45328;
	#10 counter$count = 45329;
	#10 counter$count = 45330;
	#10 counter$count = 45331;
	#10 counter$count = 45332;
	#10 counter$count = 45333;
	#10 counter$count = 45334;
	#10 counter$count = 45335;
	#10 counter$count = 45336;
	#10 counter$count = 45337;
	#10 counter$count = 45338;
	#10 counter$count = 45339;
	#10 counter$count = 45340;
	#10 counter$count = 45341;
	#10 counter$count = 45342;
	#10 counter$count = 45343;
	#10 counter$count = 45344;
	#10 counter$count = 45345;
	#10 counter$count = 45346;
	#10 counter$count = 45347;
	#10 counter$count = 45348;
	#10 counter$count = 45349;
	#10 counter$count = 45350;
	#10 counter$count = 45351;
	#10 counter$count = 45352;
	#10 counter$count = 45353;
	#10 counter$count = 45354;
	#10 counter$count = 45355;
	#10 counter$count = 45356;
	#10 counter$count = 45357;
	#10 counter$count = 45358;
	#10 counter$count = 45359;
	#10 counter$count = 45360;
	#10 counter$count = 45361;
	#10 counter$count = 45362;
	#10 counter$count = 45363;
	#10 counter$count = 45364;
	#10 counter$count = 45365;
	#10 counter$count = 45366;
	#10 counter$count = 45367;
	#10 counter$count = 45368;
	#10 counter$count = 45369;
	#10 counter$count = 45370;
	#10 counter$count = 45371;
	#10 counter$count = 45372;
	#10 counter$count = 45373;
	#10 counter$count = 45374;
	#10 counter$count = 45375;
	#10 counter$count = 45376;
	#10 counter$count = 45377;
	#10 counter$count = 45378;
	#10 counter$count = 45379;
	#10 counter$count = 45380;
	#10 counter$count = 45381;
	#10 counter$count = 45382;
	#10 counter$count = 45383;
	#10 counter$count = 45384;
	#10 counter$count = 45385;
	#10 counter$count = 45386;
	#10 counter$count = 45387;
	#10 counter$count = 45388;
	#10 counter$count = 45389;
	#10 counter$count = 45390;
	#10 counter$count = 45391;
	#10 counter$count = 45392;
	#10 counter$count = 45393;
	#10 counter$count = 45394;
	#10 counter$count = 45395;
	#10 counter$count = 45396;
	#10 counter$count = 45397;
	#10 counter$count = 45398;
	#10 counter$count = 45399;
	#10 counter$count = 45400;
	#10 counter$count = 45401;
	#10 counter$count = 45402;
	#10 counter$count = 45403;
	#10 counter$count = 45404;
	#10 counter$count = 45405;
	#10 counter$count = 45406;
	#10 counter$count = 45407;
	#10 counter$count = 45408;
	#10 counter$count = 45409;
	#10 counter$count = 45410;
	#10 counter$count = 45411;
	#10 counter$count = 45412;
	#10 counter$count = 45413;
	#10 counter$count = 45414;
	#10 counter$count = 45415;
	#10 counter$count = 45416;
	#10 counter$count = 45417;
	#10 counter$count = 45418;
	#10 counter$count = 45419;
	#10 counter$count = 45420;
	#10 counter$count = 45421;
	#10 counter$count = 45422;
	#10 counter$count = 45423;
	#10 counter$count = 45424;
	#10 counter$count = 45425;
	#10 counter$count = 45426;
	#10 counter$count = 45427;
	#10 counter$count = 45428;
	#10 counter$count = 45429;
	#10 counter$count = 45430;
	#10 counter$count = 45431;
	#10 counter$count = 45432;
	#10 counter$count = 45433;
	#10 counter$count = 45434;
	#10 counter$count = 45435;
	#10 counter$count = 45436;
	#10 counter$count = 45437;
	#10 counter$count = 45438;
	#10 counter$count = 45439;
	#10 counter$count = 45440;
	#10 counter$count = 45441;
	#10 counter$count = 45442;
	#10 counter$count = 45443;
	#10 counter$count = 45444;
	#10 counter$count = 45445;
	#10 counter$count = 45446;
	#10 counter$count = 45447;
	#10 counter$count = 45448;
	#10 counter$count = 45449;
	#10 counter$count = 45450;
	#10 counter$count = 45451;
	#10 counter$count = 45452;
	#10 counter$count = 45453;
	#10 counter$count = 45454;
	#10 counter$count = 45455;
	#10 counter$count = 45456;
	#10 counter$count = 45457;
	#10 counter$count = 45458;
	#10 counter$count = 45459;
	#10 counter$count = 45460;
	#10 counter$count = 45461;
	#10 counter$count = 45462;
	#10 counter$count = 45463;
	#10 counter$count = 45464;
	#10 counter$count = 45465;
	#10 counter$count = 45466;
	#10 counter$count = 45467;
	#10 counter$count = 45468;
	#10 counter$count = 45469;
	#10 counter$count = 45470;
	#10 counter$count = 45471;
	#10 counter$count = 45472;
	#10 counter$count = 45473;
	#10 counter$count = 45474;
	#10 counter$count = 45475;
	#10 counter$count = 45476;
	#10 counter$count = 45477;
	#10 counter$count = 45478;
	#10 counter$count = 45479;
	#10 counter$count = 45480;
	#10 counter$count = 45481;
	#10 counter$count = 45482;
	#10 counter$count = 45483;
	#10 counter$count = 45484;
	#10 counter$count = 45485;
	#10 counter$count = 45486;
	#10 counter$count = 45487;
	#10 counter$count = 45488;
	#10 counter$count = 45489;
	#10 counter$count = 45490;
	#10 counter$count = 45491;
	#10 counter$count = 45492;
	#10 counter$count = 45493;
	#10 counter$count = 45494;
	#10 counter$count = 45495;
	#10 counter$count = 45496;
	#10 counter$count = 45497;
	#10 counter$count = 45498;
	#10 counter$count = 45499;
	#10 counter$count = 45500;
	#10 counter$count = 45501;
	#10 counter$count = 45502;
	#10 counter$count = 45503;
	#10 counter$count = 45504;
	#10 counter$count = 45505;
	#10 counter$count = 45506;
	#10 counter$count = 45507;
	#10 counter$count = 45508;
	#10 counter$count = 45509;
	#10 counter$count = 45510;
	#10 counter$count = 45511;
	#10 counter$count = 45512;
	#10 counter$count = 45513;
	#10 counter$count = 45514;
	#10 counter$count = 45515;
	#10 counter$count = 45516;
	#10 counter$count = 45517;
	#10 counter$count = 45518;
	#10 counter$count = 45519;
	#10 counter$count = 45520;
	#10 counter$count = 45521;
	#10 counter$count = 45522;
	#10 counter$count = 45523;
	#10 counter$count = 45524;
	#10 counter$count = 45525;
	#10 counter$count = 45526;
	#10 counter$count = 45527;
	#10 counter$count = 45528;
	#10 counter$count = 45529;
	#10 counter$count = 45530;
	#10 counter$count = 45531;
	#10 counter$count = 45532;
	#10 counter$count = 45533;
	#10 counter$count = 45534;
	#10 counter$count = 45535;
	#10 counter$count = 45536;
	#10 counter$count = 45537;
	#10 counter$count = 45538;
	#10 counter$count = 45539;
	#10 counter$count = 45540;
	#10 counter$count = 45541;
	#10 counter$count = 45542;
	#10 counter$count = 45543;
	#10 counter$count = 45544;
	#10 counter$count = 45545;
	#10 counter$count = 45546;
	#10 counter$count = 45547;
	#10 counter$count = 45548;
	#10 counter$count = 45549;
	#10 counter$count = 45550;
	#10 counter$count = 45551;
	#10 counter$count = 45552;
	#10 counter$count = 45553;
	#10 counter$count = 45554;
	#10 counter$count = 45555;
	#10 counter$count = 45556;
	#10 counter$count = 45557;
	#10 counter$count = 45558;
	#10 counter$count = 45559;
	#10 counter$count = 45560;
	#10 counter$count = 45561;
	#10 counter$count = 45562;
	#10 counter$count = 45563;
	#10 counter$count = 45564;
	#10 counter$count = 45565;
	#10 counter$count = 45566;
	#10 counter$count = 45567;
	#10 counter$count = 45568;
	#10 counter$count = 45569;
	#10 counter$count = 45570;
	#10 counter$count = 45571;
	#10 counter$count = 45572;
	#10 counter$count = 45573;
	#10 counter$count = 45574;
	#10 counter$count = 45575;
	#10 counter$count = 45576;
	#10 counter$count = 45577;
	#10 counter$count = 45578;
	#10 counter$count = 45579;
	#10 counter$count = 45580;
	#10 counter$count = 45581;
	#10 counter$count = 45582;
	#10 counter$count = 45583;
	#10 counter$count = 45584;
	#10 counter$count = 45585;
	#10 counter$count = 45586;
	#10 counter$count = 45587;
	#10 counter$count = 45588;
	#10 counter$count = 45589;
	#10 counter$count = 45590;
	#10 counter$count = 45591;
	#10 counter$count = 45592;
	#10 counter$count = 45593;
	#10 counter$count = 45594;
	#10 counter$count = 45595;
	#10 counter$count = 45596;
	#10 counter$count = 45597;
	#10 counter$count = 45598;
	#10 counter$count = 45599;
	#10 counter$count = 45600;
	#10 counter$count = 45601;
	#10 counter$count = 45602;
	#10 counter$count = 45603;
	#10 counter$count = 45604;
	#10 counter$count = 45605;
	#10 counter$count = 45606;
	#10 counter$count = 45607;
	#10 counter$count = 45608;
	#10 counter$count = 45609;
	#10 counter$count = 45610;
	#10 counter$count = 45611;
	#10 counter$count = 45612;
	#10 counter$count = 45613;
	#10 counter$count = 45614;
	#10 counter$count = 45615;
	#10 counter$count = 45616;
	#10 counter$count = 45617;
	#10 counter$count = 45618;
	#10 counter$count = 45619;
	#10 counter$count = 45620;
	#10 counter$count = 45621;
	#10 counter$count = 45622;
	#10 counter$count = 45623;
	#10 counter$count = 45624;
	#10 counter$count = 45625;
	#10 counter$count = 45626;
	#10 counter$count = 45627;
	#10 counter$count = 45628;
	#10 counter$count = 45629;
	#10 counter$count = 45630;
	#10 counter$count = 45631;
	#10 counter$count = 45632;
	#10 counter$count = 45633;
	#10 counter$count = 45634;
	#10 counter$count = 45635;
	#10 counter$count = 45636;
	#10 counter$count = 45637;
	#10 counter$count = 45638;
	#10 counter$count = 45639;
	#10 counter$count = 45640;
	#10 counter$count = 45641;
	#10 counter$count = 45642;
	#10 counter$count = 45643;
	#10 counter$count = 45644;
	#10 counter$count = 45645;
	#10 counter$count = 45646;
	#10 counter$count = 45647;
	#10 counter$count = 45648;
	#10 counter$count = 45649;
	#10 counter$count = 45650;
	#10 counter$count = 45651;
	#10 counter$count = 45652;
	#10 counter$count = 45653;
	#10 counter$count = 45654;
	#10 counter$count = 45655;
	#10 counter$count = 45656;
	#10 counter$count = 45657;
	#10 counter$count = 45658;
	#10 counter$count = 45659;
	#10 counter$count = 45660;
	#10 counter$count = 45661;
	#10 counter$count = 45662;
	#10 counter$count = 45663;
	#10 counter$count = 45664;
	#10 counter$count = 45665;
	#10 counter$count = 45666;
	#10 counter$count = 45667;
	#10 counter$count = 45668;
	#10 counter$count = 45669;
	#10 counter$count = 45670;
	#10 counter$count = 45671;
	#10 counter$count = 45672;
	#10 counter$count = 45673;
	#10 counter$count = 45674;
	#10 counter$count = 45675;
	#10 counter$count = 45676;
	#10 counter$count = 45677;
	#10 counter$count = 45678;
	#10 counter$count = 45679;
	#10 counter$count = 45680;
	#10 counter$count = 45681;
	#10 counter$count = 45682;
	#10 counter$count = 45683;
	#10 counter$count = 45684;
	#10 counter$count = 45685;
	#10 counter$count = 45686;
	#10 counter$count = 45687;
	#10 counter$count = 45688;
	#10 counter$count = 45689;
	#10 counter$count = 45690;
	#10 counter$count = 45691;
	#10 counter$count = 45692;
	#10 counter$count = 45693;
	#10 counter$count = 45694;
	#10 counter$count = 45695;
	#10 counter$count = 45696;
	#10 counter$count = 45697;
	#10 counter$count = 45698;
	#10 counter$count = 45699;
	#10 counter$count = 45700;
	#10 counter$count = 45701;
	#10 counter$count = 45702;
	#10 counter$count = 45703;
	#10 counter$count = 45704;
	#10 counter$count = 45705;
	#10 counter$count = 45706;
	#10 counter$count = 45707;
	#10 counter$count = 45708;
	#10 counter$count = 45709;
	#10 counter$count = 45710;
	#10 counter$count = 45711;
	#10 counter$count = 45712;
	#10 counter$count = 45713;
	#10 counter$count = 45714;
	#10 counter$count = 45715;
	#10 counter$count = 45716;
	#10 counter$count = 45717;
	#10 counter$count = 45718;
	#10 counter$count = 45719;
	#10 counter$count = 45720;
	#10 counter$count = 45721;
	#10 counter$count = 45722;
	#10 counter$count = 45723;
	#10 counter$count = 45724;
	#10 counter$count = 45725;
	#10 counter$count = 45726;
	#10 counter$count = 45727;
	#10 counter$count = 45728;
	#10 counter$count = 45729;
	#10 counter$count = 45730;
	#10 counter$count = 45731;
	#10 counter$count = 45732;
	#10 counter$count = 45733;
	#10 counter$count = 45734;
	#10 counter$count = 45735;
	#10 counter$count = 45736;
	#10 counter$count = 45737;
	#10 counter$count = 45738;
	#10 counter$count = 45739;
	#10 counter$count = 45740;
	#10 counter$count = 45741;
	#10 counter$count = 45742;
	#10 counter$count = 45743;
	#10 counter$count = 45744;
	#10 counter$count = 45745;
	#10 counter$count = 45746;
	#10 counter$count = 45747;
	#10 counter$count = 45748;
	#10 counter$count = 45749;
	#10 counter$count = 45750;
	#10 counter$count = 45751;
	#10 counter$count = 45752;
	#10 counter$count = 45753;
	#10 counter$count = 45754;
	#10 counter$count = 45755;
	#10 counter$count = 45756;
	#10 counter$count = 45757;
	#10 counter$count = 45758;
	#10 counter$count = 45759;
	#10 counter$count = 45760;
	#10 counter$count = 45761;
	#10 counter$count = 45762;
	#10 counter$count = 45763;
	#10 counter$count = 45764;
	#10 counter$count = 45765;
	#10 counter$count = 45766;
	#10 counter$count = 45767;
	#10 counter$count = 45768;
	#10 counter$count = 45769;
	#10 counter$count = 45770;
	#10 counter$count = 45771;
	#10 counter$count = 45772;
	#10 counter$count = 45773;
	#10 counter$count = 45774;
	#10 counter$count = 45775;
	#10 counter$count = 45776;
	#10 counter$count = 45777;
	#10 counter$count = 45778;
	#10 counter$count = 45779;
	#10 counter$count = 45780;
	#10 counter$count = 45781;
	#10 counter$count = 45782;
	#10 counter$count = 45783;
	#10 counter$count = 45784;
	#10 counter$count = 45785;
	#10 counter$count = 45786;
	#10 counter$count = 45787;
	#10 counter$count = 45788;
	#10 counter$count = 45789;
	#10 counter$count = 45790;
	#10 counter$count = 45791;
	#10 counter$count = 45792;
	#10 counter$count = 45793;
	#10 counter$count = 45794;
	#10 counter$count = 45795;
	#10 counter$count = 45796;
	#10 counter$count = 45797;
	#10 counter$count = 45798;
	#10 counter$count = 45799;
	#10 counter$count = 45800;
	#10 counter$count = 45801;
	#10 counter$count = 45802;
	#10 counter$count = 45803;
	#10 counter$count = 45804;
	#10 counter$count = 45805;
	#10 counter$count = 45806;
	#10 counter$count = 45807;
	#10 counter$count = 45808;
	#10 counter$count = 45809;
	#10 counter$count = 45810;
	#10 counter$count = 45811;
	#10 counter$count = 45812;
	#10 counter$count = 45813;
	#10 counter$count = 45814;
	#10 counter$count = 45815;
	#10 counter$count = 45816;
	#10 counter$count = 45817;
	#10 counter$count = 45818;
	#10 counter$count = 45819;
	#10 counter$count = 45820;
	#10 counter$count = 45821;
	#10 counter$count = 45822;
	#10 counter$count = 45823;
	#10 counter$count = 45824;
	#10 counter$count = 45825;
	#10 counter$count = 45826;
	#10 counter$count = 45827;
	#10 counter$count = 45828;
	#10 counter$count = 45829;
	#10 counter$count = 45830;
	#10 counter$count = 45831;
	#10 counter$count = 45832;
	#10 counter$count = 45833;
	#10 counter$count = 45834;
	#10 counter$count = 45835;
	#10 counter$count = 45836;
	#10 counter$count = 45837;
	#10 counter$count = 45838;
	#10 counter$count = 45839;
	#10 counter$count = 45840;
	#10 counter$count = 45841;
	#10 counter$count = 45842;
	#10 counter$count = 45843;
	#10 counter$count = 45844;
	#10 counter$count = 45845;
	#10 counter$count = 45846;
	#10 counter$count = 45847;
	#10 counter$count = 45848;
	#10 counter$count = 45849;
	#10 counter$count = 45850;
	#10 counter$count = 45851;
	#10 counter$count = 45852;
	#10 counter$count = 45853;
	#10 counter$count = 45854;
	#10 counter$count = 45855;
	#10 counter$count = 45856;
	#10 counter$count = 45857;
	#10 counter$count = 45858;
	#10 counter$count = 45859;
	#10 counter$count = 45860;
	#10 counter$count = 45861;
	#10 counter$count = 45862;
	#10 counter$count = 45863;
	#10 counter$count = 45864;
	#10 counter$count = 45865;
	#10 counter$count = 45866;
	#10 counter$count = 45867;
	#10 counter$count = 45868;
	#10 counter$count = 45869;
	#10 counter$count = 45870;
	#10 counter$count = 45871;
	#10 counter$count = 45872;
	#10 counter$count = 45873;
	#10 counter$count = 45874;
	#10 counter$count = 45875;
	#10 counter$count = 45876;
	#10 counter$count = 45877;
	#10 counter$count = 45878;
	#10 counter$count = 45879;
	#10 counter$count = 45880;
	#10 counter$count = 45881;
	#10 counter$count = 45882;
	#10 counter$count = 45883;
	#10 counter$count = 45884;
	#10 counter$count = 45885;
	#10 counter$count = 45886;
	#10 counter$count = 45887;
	#10 counter$count = 45888;
	#10 counter$count = 45889;
	#10 counter$count = 45890;
	#10 counter$count = 45891;
	#10 counter$count = 45892;
	#10 counter$count = 45893;
	#10 counter$count = 45894;
	#10 counter$count = 45895;
	#10 counter$count = 45896;
	#10 counter$count = 45897;
	#10 counter$count = 45898;
	#10 counter$count = 45899;
	#10 counter$count = 45900;
	#10 counter$count = 45901;
	#10 counter$count = 45902;
	#10 counter$count = 45903;
	#10 counter$count = 45904;
	#10 counter$count = 45905;
	#10 counter$count = 45906;
	#10 counter$count = 45907;
	#10 counter$count = 45908;
	#10 counter$count = 45909;
	#10 counter$count = 45910;
	#10 counter$count = 45911;
	#10 counter$count = 45912;
	#10 counter$count = 45913;
	#10 counter$count = 45914;
	#10 counter$count = 45915;
	#10 counter$count = 45916;
	#10 counter$count = 45917;
	#10 counter$count = 45918;
	#10 counter$count = 45919;
	#10 counter$count = 45920;
	#10 counter$count = 45921;
	#10 counter$count = 45922;
	#10 counter$count = 45923;
	#10 counter$count = 45924;
	#10 counter$count = 45925;
	#10 counter$count = 45926;
	#10 counter$count = 45927;
	#10 counter$count = 45928;
	#10 counter$count = 45929;
	#10 counter$count = 45930;
	#10 counter$count = 45931;
	#10 counter$count = 45932;
	#10 counter$count = 45933;
	#10 counter$count = 45934;
	#10 counter$count = 45935;
	#10 counter$count = 45936;
	#10 counter$count = 45937;
	#10 counter$count = 45938;
	#10 counter$count = 45939;
	#10 counter$count = 45940;
	#10 counter$count = 45941;
	#10 counter$count = 45942;
	#10 counter$count = 45943;
	#10 counter$count = 45944;
	#10 counter$count = 45945;
	#10 counter$count = 45946;
	#10 counter$count = 45947;
	#10 counter$count = 45948;
	#10 counter$count = 45949;
	#10 counter$count = 45950;
	#10 counter$count = 45951;
	#10 counter$count = 45952;
	#10 counter$count = 45953;
	#10 counter$count = 45954;
	#10 counter$count = 45955;
	#10 counter$count = 45956;
	#10 counter$count = 45957;
	#10 counter$count = 45958;
	#10 counter$count = 45959;
	#10 counter$count = 45960;
	#10 counter$count = 45961;
	#10 counter$count = 45962;
	#10 counter$count = 45963;
	#10 counter$count = 45964;
	#10 counter$count = 45965;
	#10 counter$count = 45966;
	#10 counter$count = 45967;
	#10 counter$count = 45968;
	#10 counter$count = 45969;
	#10 counter$count = 45970;
	#10 counter$count = 45971;
	#10 counter$count = 45972;
	#10 counter$count = 45973;
	#10 counter$count = 45974;
	#10 counter$count = 45975;
	#10 counter$count = 45976;
	#10 counter$count = 45977;
	#10 counter$count = 45978;
	#10 counter$count = 45979;
	#10 counter$count = 45980;
	#10 counter$count = 45981;
	#10 counter$count = 45982;
	#10 counter$count = 45983;
	#10 counter$count = 45984;
	#10 counter$count = 45985;
	#10 counter$count = 45986;
	#10 counter$count = 45987;
	#10 counter$count = 45988;
	#10 counter$count = 45989;
	#10 counter$count = 45990;
	#10 counter$count = 45991;
	#10 counter$count = 45992;
	#10 counter$count = 45993;
	#10 counter$count = 45994;
	#10 counter$count = 45995;
	#10 counter$count = 45996;
	#10 counter$count = 45997;
	#10 counter$count = 45998;
	#10 counter$count = 45999;
	#10 counter$count = 46000;
	#10 counter$count = 46001;
	#10 counter$count = 46002;
	#10 counter$count = 46003;
	#10 counter$count = 46004;
	#10 counter$count = 46005;
	#10 counter$count = 46006;
	#10 counter$count = 46007;
	#10 counter$count = 46008;
	#10 counter$count = 46009;
	#10 counter$count = 46010;
	#10 counter$count = 46011;
	#10 counter$count = 46012;
	#10 counter$count = 46013;
	#10 counter$count = 46014;
	#10 counter$count = 46015;
	#10 counter$count = 46016;
	#10 counter$count = 46017;
	#10 counter$count = 46018;
	#10 counter$count = 46019;
	#10 counter$count = 46020;
	#10 counter$count = 46021;
	#10 counter$count = 46022;
	#10 counter$count = 46023;
	#10 counter$count = 46024;
	#10 counter$count = 46025;
	#10 counter$count = 46026;
	#10 counter$count = 46027;
	#10 counter$count = 46028;
	#10 counter$count = 46029;
	#10 counter$count = 46030;
	#10 counter$count = 46031;
	#10 counter$count = 46032;
	#10 counter$count = 46033;
	#10 counter$count = 46034;
	#10 counter$count = 46035;
	#10 counter$count = 46036;
	#10 counter$count = 46037;
	#10 counter$count = 46038;
	#10 counter$count = 46039;
	#10 counter$count = 46040;
	#10 counter$count = 46041;
	#10 counter$count = 46042;
	#10 counter$count = 46043;
	#10 counter$count = 46044;
	#10 counter$count = 46045;
	#10 counter$count = 46046;
	#10 counter$count = 46047;
	#10 counter$count = 46048;
	#10 counter$count = 46049;
	#10 counter$count = 46050;
	#10 counter$count = 46051;
	#10 counter$count = 46052;
	#10 counter$count = 46053;
	#10 counter$count = 46054;
	#10 counter$count = 46055;
	#10 counter$count = 46056;
	#10 counter$count = 46057;
	#10 counter$count = 46058;
	#10 counter$count = 46059;
	#10 counter$count = 46060;
	#10 counter$count = 46061;
	#10 counter$count = 46062;
	#10 counter$count = 46063;
	#10 counter$count = 46064;
	#10 counter$count = 46065;
	#10 counter$count = 46066;
	#10 counter$count = 46067;
	#10 counter$count = 46068;
	#10 counter$count = 46069;
	#10 counter$count = 46070;
	#10 counter$count = 46071;
	#10 counter$count = 46072;
	#10 counter$count = 46073;
	#10 counter$count = 46074;
	#10 counter$count = 46075;
	#10 counter$count = 46076;
	#10 counter$count = 46077;
	#10 counter$count = 46078;
	#10 counter$count = 46079;
	#10 counter$count = 46080;
	#10 counter$count = 46081;
	#10 counter$count = 46082;
	#10 counter$count = 46083;
	#10 counter$count = 46084;
	#10 counter$count = 46085;
	#10 counter$count = 46086;
	#10 counter$count = 46087;
	#10 counter$count = 46088;
	#10 counter$count = 46089;
	#10 counter$count = 46090;
	#10 counter$count = 46091;
	#10 counter$count = 46092;
	#10 counter$count = 46093;
	#10 counter$count = 46094;
	#10 counter$count = 46095;
	#10 counter$count = 46096;
	#10 counter$count = 46097;
	#10 counter$count = 46098;
	#10 counter$count = 46099;
	#10 counter$count = 46100;
	#10 counter$count = 46101;
	#10 counter$count = 46102;
	#10 counter$count = 46103;
	#10 counter$count = 46104;
	#10 counter$count = 46105;
	#10 counter$count = 46106;
	#10 counter$count = 46107;
	#10 counter$count = 46108;
	#10 counter$count = 46109;
	#10 counter$count = 46110;
	#10 counter$count = 46111;
	#10 counter$count = 46112;
	#10 counter$count = 46113;
	#10 counter$count = 46114;
	#10 counter$count = 46115;
	#10 counter$count = 46116;
	#10 counter$count = 46117;
	#10 counter$count = 46118;
	#10 counter$count = 46119;
	#10 counter$count = 46120;
	#10 counter$count = 46121;
	#10 counter$count = 46122;
	#10 counter$count = 46123;
	#10 counter$count = 46124;
	#10 counter$count = 46125;
	#10 counter$count = 46126;
	#10 counter$count = 46127;
	#10 counter$count = 46128;
	#10 counter$count = 46129;
	#10 counter$count = 46130;
	#10 counter$count = 46131;
	#10 counter$count = 46132;
	#10 counter$count = 46133;
	#10 counter$count = 46134;
	#10 counter$count = 46135;
	#10 counter$count = 46136;
	#10 counter$count = 46137;
	#10 counter$count = 46138;
	#10 counter$count = 46139;
	#10 counter$count = 46140;
	#10 counter$count = 46141;
	#10 counter$count = 46142;
	#10 counter$count = 46143;
	#10 counter$count = 46144;
	#10 counter$count = 46145;
	#10 counter$count = 46146;
	#10 counter$count = 46147;
	#10 counter$count = 46148;
	#10 counter$count = 46149;
	#10 counter$count = 46150;
	#10 counter$count = 46151;
	#10 counter$count = 46152;
	#10 counter$count = 46153;
	#10 counter$count = 46154;
	#10 counter$count = 46155;
	#10 counter$count = 46156;
	#10 counter$count = 46157;
	#10 counter$count = 46158;
	#10 counter$count = 46159;
	#10 counter$count = 46160;
	#10 counter$count = 46161;
	#10 counter$count = 46162;
	#10 counter$count = 46163;
	#10 counter$count = 46164;
	#10 counter$count = 46165;
	#10 counter$count = 46166;
	#10 counter$count = 46167;
	#10 counter$count = 46168;
	#10 counter$count = 46169;
	#10 counter$count = 46170;
	#10 counter$count = 46171;
	#10 counter$count = 46172;
	#10 counter$count = 46173;
	#10 counter$count = 46174;
	#10 counter$count = 46175;
	#10 counter$count = 46176;
	#10 counter$count = 46177;
	#10 counter$count = 46178;
	#10 counter$count = 46179;
	#10 counter$count = 46180;
	#10 counter$count = 46181;
	#10 counter$count = 46182;
	#10 counter$count = 46183;
	#10 counter$count = 46184;
	#10 counter$count = 46185;
	#10 counter$count = 46186;
	#10 counter$count = 46187;
	#10 counter$count = 46188;
	#10 counter$count = 46189;
	#10 counter$count = 46190;
	#10 counter$count = 46191;
	#10 counter$count = 46192;
	#10 counter$count = 46193;
	#10 counter$count = 46194;
	#10 counter$count = 46195;
	#10 counter$count = 46196;
	#10 counter$count = 46197;
	#10 counter$count = 46198;
	#10 counter$count = 46199;
	#10 counter$count = 46200;
	#10 counter$count = 46201;
	#10 counter$count = 46202;
	#10 counter$count = 46203;
	#10 counter$count = 46204;
	#10 counter$count = 46205;
	#10 counter$count = 46206;
	#10 counter$count = 46207;
	#10 counter$count = 46208;
	#10 counter$count = 46209;
	#10 counter$count = 46210;
	#10 counter$count = 46211;
	#10 counter$count = 46212;
	#10 counter$count = 46213;
	#10 counter$count = 46214;
	#10 counter$count = 46215;
	#10 counter$count = 46216;
	#10 counter$count = 46217;
	#10 counter$count = 46218;
	#10 counter$count = 46219;
	#10 counter$count = 46220;
	#10 counter$count = 46221;
	#10 counter$count = 46222;
	#10 counter$count = 46223;
	#10 counter$count = 46224;
	#10 counter$count = 46225;
	#10 counter$count = 46226;
	#10 counter$count = 46227;
	#10 counter$count = 46228;
	#10 counter$count = 46229;
	#10 counter$count = 46230;
	#10 counter$count = 46231;
	#10 counter$count = 46232;
	#10 counter$count = 46233;
	#10 counter$count = 46234;
	#10 counter$count = 46235;
	#10 counter$count = 46236;
	#10 counter$count = 46237;
	#10 counter$count = 46238;
	#10 counter$count = 46239;
	#10 counter$count = 46240;
	#10 counter$count = 46241;
	#10 counter$count = 46242;
	#10 counter$count = 46243;
	#10 counter$count = 46244;
	#10 counter$count = 46245;
	#10 counter$count = 46246;
	#10 counter$count = 46247;
	#10 counter$count = 46248;
	#10 counter$count = 46249;
	#10 counter$count = 46250;
	#10 counter$count = 46251;
	#10 counter$count = 46252;
	#10 counter$count = 46253;
	#10 counter$count = 46254;
	#10 counter$count = 46255;
	#10 counter$count = 46256;
	#10 counter$count = 46257;
	#10 counter$count = 46258;
	#10 counter$count = 46259;
	#10 counter$count = 46260;
	#10 counter$count = 46261;
	#10 counter$count = 46262;
	#10 counter$count = 46263;
	#10 counter$count = 46264;
	#10 counter$count = 46265;
	#10 counter$count = 46266;
	#10 counter$count = 46267;
	#10 counter$count = 46268;
	#10 counter$count = 46269;
	#10 counter$count = 46270;
	#10 counter$count = 46271;
	#10 counter$count = 46272;
	#10 counter$count = 46273;
	#10 counter$count = 46274;
	#10 counter$count = 46275;
	#10 counter$count = 46276;
	#10 counter$count = 46277;
	#10 counter$count = 46278;
	#10 counter$count = 46279;
	#10 counter$count = 46280;
	#10 counter$count = 46281;
	#10 counter$count = 46282;
	#10 counter$count = 46283;
	#10 counter$count = 46284;
	#10 counter$count = 46285;
	#10 counter$count = 46286;
	#10 counter$count = 46287;
	#10 counter$count = 46288;
	#10 counter$count = 46289;
	#10 counter$count = 46290;
	#10 counter$count = 46291;
	#10 counter$count = 46292;
	#10 counter$count = 46293;
	#10 counter$count = 46294;
	#10 counter$count = 46295;
	#10 counter$count = 46296;
	#10 counter$count = 46297;
	#10 counter$count = 46298;
	#10 counter$count = 46299;
	#10 counter$count = 46300;
	#10 counter$count = 46301;
	#10 counter$count = 46302;
	#10 counter$count = 46303;
	#10 counter$count = 46304;
	#10 counter$count = 46305;
	#10 counter$count = 46306;
	#10 counter$count = 46307;
	#10 counter$count = 46308;
	#10 counter$count = 46309;
	#10 counter$count = 46310;
	#10 counter$count = 46311;
	#10 counter$count = 46312;
	#10 counter$count = 46313;
	#10 counter$count = 46314;
	#10 counter$count = 46315;
	#10 counter$count = 46316;
	#10 counter$count = 46317;
	#10 counter$count = 46318;
	#10 counter$count = 46319;
	#10 counter$count = 46320;
	#10 counter$count = 46321;
	#10 counter$count = 46322;
	#10 counter$count = 46323;
	#10 counter$count = 46324;
	#10 counter$count = 46325;
	#10 counter$count = 46326;
	#10 counter$count = 46327;
	#10 counter$count = 46328;
	#10 counter$count = 46329;
	#10 counter$count = 46330;
	#10 counter$count = 46331;
	#10 counter$count = 46332;
	#10 counter$count = 46333;
	#10 counter$count = 46334;
	#10 counter$count = 46335;
	#10 counter$count = 46336;
	#10 counter$count = 46337;
	#10 counter$count = 46338;
	#10 counter$count = 46339;
	#10 counter$count = 46340;
	#10 counter$count = 46341;
	#10 counter$count = 46342;
	#10 counter$count = 46343;
	#10 counter$count = 46344;
	#10 counter$count = 46345;
	#10 counter$count = 46346;
	#10 counter$count = 46347;
	#10 counter$count = 46348;
	#10 counter$count = 46349;
	#10 counter$count = 46350;
	#10 counter$count = 46351;
	#10 counter$count = 46352;
	#10 counter$count = 46353;
	#10 counter$count = 46354;
	#10 counter$count = 46355;
	#10 counter$count = 46356;
	#10 counter$count = 46357;
	#10 counter$count = 46358;
	#10 counter$count = 46359;
	#10 counter$count = 46360;
	#10 counter$count = 46361;
	#10 counter$count = 46362;
	#10 counter$count = 46363;
	#10 counter$count = 46364;
	#10 counter$count = 46365;
	#10 counter$count = 46366;
	#10 counter$count = 46367;
	#10 counter$count = 46368;
	#10 counter$count = 46369;
	#10 counter$count = 46370;
	#10 counter$count = 46371;
	#10 counter$count = 46372;
	#10 counter$count = 46373;
	#10 counter$count = 46374;
	#10 counter$count = 46375;
	#10 counter$count = 46376;
	#10 counter$count = 46377;
	#10 counter$count = 46378;
	#10 counter$count = 46379;
	#10 counter$count = 46380;
	#10 counter$count = 46381;
	#10 counter$count = 46382;
	#10 counter$count = 46383;
	#10 counter$count = 46384;
	#10 counter$count = 46385;
	#10 counter$count = 46386;
	#10 counter$count = 46387;
	#10 counter$count = 46388;
	#10 counter$count = 46389;
	#10 counter$count = 46390;
	#10 counter$count = 46391;
	#10 counter$count = 46392;
	#10 counter$count = 46393;
	#10 counter$count = 46394;
	#10 counter$count = 46395;
	#10 counter$count = 46396;
	#10 counter$count = 46397;
	#10 counter$count = 46398;
	#10 counter$count = 46399;
	#10 counter$count = 46400;
	#10 counter$count = 46401;
	#10 counter$count = 46402;
	#10 counter$count = 46403;
	#10 counter$count = 46404;
	#10 counter$count = 46405;
	#10 counter$count = 46406;
	#10 counter$count = 46407;
	#10 counter$count = 46408;
	#10 counter$count = 46409;
	#10 counter$count = 46410;
	#10 counter$count = 46411;
	#10 counter$count = 46412;
	#10 counter$count = 46413;
	#10 counter$count = 46414;
	#10 counter$count = 46415;
	#10 counter$count = 46416;
	#10 counter$count = 46417;
	#10 counter$count = 46418;
	#10 counter$count = 46419;
	#10 counter$count = 46420;
	#10 counter$count = 46421;
	#10 counter$count = 46422;
	#10 counter$count = 46423;
	#10 counter$count = 46424;
	#10 counter$count = 46425;
	#10 counter$count = 46426;
	#10 counter$count = 46427;
	#10 counter$count = 46428;
	#10 counter$count = 46429;
	#10 counter$count = 46430;
	#10 counter$count = 46431;
	#10 counter$count = 46432;
	#10 counter$count = 46433;
	#10 counter$count = 46434;
	#10 counter$count = 46435;
	#10 counter$count = 46436;
	#10 counter$count = 46437;
	#10 counter$count = 46438;
	#10 counter$count = 46439;
	#10 counter$count = 46440;
	#10 counter$count = 46441;
	#10 counter$count = 46442;
	#10 counter$count = 46443;
	#10 counter$count = 46444;
	#10 counter$count = 46445;
	#10 counter$count = 46446;
	#10 counter$count = 46447;
	#10 counter$count = 46448;
	#10 counter$count = 46449;
	#10 counter$count = 46450;
	#10 counter$count = 46451;
	#10 counter$count = 46452;
	#10 counter$count = 46453;
	#10 counter$count = 46454;
	#10 counter$count = 46455;
	#10 counter$count = 46456;
	#10 counter$count = 46457;
	#10 counter$count = 46458;
	#10 counter$count = 46459;
	#10 counter$count = 46460;
	#10 counter$count = 46461;
	#10 counter$count = 46462;
	#10 counter$count = 46463;
	#10 counter$count = 46464;
	#10 counter$count = 46465;
	#10 counter$count = 46466;
	#10 counter$count = 46467;
	#10 counter$count = 46468;
	#10 counter$count = 46469;
	#10 counter$count = 46470;
	#10 counter$count = 46471;
	#10 counter$count = 46472;
	#10 counter$count = 46473;
	#10 counter$count = 46474;
	#10 counter$count = 46475;
	#10 counter$count = 46476;
	#10 counter$count = 46477;
	#10 counter$count = 46478;
	#10 counter$count = 46479;
	#10 counter$count = 46480;
	#10 counter$count = 46481;
	#10 counter$count = 46482;
	#10 counter$count = 46483;
	#10 counter$count = 46484;
	#10 counter$count = 46485;
	#10 counter$count = 46486;
	#10 counter$count = 46487;
	#10 counter$count = 46488;
	#10 counter$count = 46489;
	#10 counter$count = 46490;
	#10 counter$count = 46491;
	#10 counter$count = 46492;
	#10 counter$count = 46493;
	#10 counter$count = 46494;
	#10 counter$count = 46495;
	#10 counter$count = 46496;
	#10 counter$count = 46497;
	#10 counter$count = 46498;
	#10 counter$count = 46499;
	#10 counter$count = 46500;
	#10 counter$count = 46501;
	#10 counter$count = 46502;
	#10 counter$count = 46503;
	#10 counter$count = 46504;
	#10 counter$count = 46505;
	#10 counter$count = 46506;
	#10 counter$count = 46507;
	#10 counter$count = 46508;
	#10 counter$count = 46509;
	#10 counter$count = 46510;
	#10 counter$count = 46511;
	#10 counter$count = 46512;
	#10 counter$count = 46513;
	#10 counter$count = 46514;
	#10 counter$count = 46515;
	#10 counter$count = 46516;
	#10 counter$count = 46517;
	#10 counter$count = 46518;
	#10 counter$count = 46519;
	#10 counter$count = 46520;
	#10 counter$count = 46521;
	#10 counter$count = 46522;
	#10 counter$count = 46523;
	#10 counter$count = 46524;
	#10 counter$count = 46525;
	#10 counter$count = 46526;
	#10 counter$count = 46527;
	#10 counter$count = 46528;
	#10 counter$count = 46529;
	#10 counter$count = 46530;
	#10 counter$count = 46531;
	#10 counter$count = 46532;
	#10 counter$count = 46533;
	#10 counter$count = 46534;
	#10 counter$count = 46535;
	#10 counter$count = 46536;
	#10 counter$count = 46537;
	#10 counter$count = 46538;
	#10 counter$count = 46539;
	#10 counter$count = 46540;
	#10 counter$count = 46541;
	#10 counter$count = 46542;
	#10 counter$count = 46543;
	#10 counter$count = 46544;
	#10 counter$count = 46545;
	#10 counter$count = 46546;
	#10 counter$count = 46547;
	#10 counter$count = 46548;
	#10 counter$count = 46549;
	#10 counter$count = 46550;
	#10 counter$count = 46551;
	#10 counter$count = 46552;
	#10 counter$count = 46553;
	#10 counter$count = 46554;
	#10 counter$count = 46555;
	#10 counter$count = 46556;
	#10 counter$count = 46557;
	#10 counter$count = 46558;
	#10 counter$count = 46559;
	#10 counter$count = 46560;
	#10 counter$count = 46561;
	#10 counter$count = 46562;
	#10 counter$count = 46563;
	#10 counter$count = 46564;
	#10 counter$count = 46565;
	#10 counter$count = 46566;
	#10 counter$count = 46567;
	#10 counter$count = 46568;
	#10 counter$count = 46569;
	#10 counter$count = 46570;
	#10 counter$count = 46571;
	#10 counter$count = 46572;
	#10 counter$count = 46573;
	#10 counter$count = 46574;
	#10 counter$count = 46575;
	#10 counter$count = 46576;
	#10 counter$count = 46577;
	#10 counter$count = 46578;
	#10 counter$count = 46579;
	#10 counter$count = 46580;
	#10 counter$count = 46581;
	#10 counter$count = 46582;
	#10 counter$count = 46583;
	#10 counter$count = 46584;
	#10 counter$count = 46585;
	#10 counter$count = 46586;
	#10 counter$count = 46587;
	#10 counter$count = 46588;
	#10 counter$count = 46589;
	#10 counter$count = 46590;
	#10 counter$count = 46591;
	#10 counter$count = 46592;
	#10 counter$count = 46593;
	#10 counter$count = 46594;
	#10 counter$count = 46595;
	#10 counter$count = 46596;
	#10 counter$count = 46597;
	#10 counter$count = 46598;
	#10 counter$count = 46599;
	#10 counter$count = 46600;
	#10 counter$count = 46601;
	#10 counter$count = 46602;
	#10 counter$count = 46603;
	#10 counter$count = 46604;
	#10 counter$count = 46605;
	#10 counter$count = 46606;
	#10 counter$count = 46607;
	#10 counter$count = 46608;
	#10 counter$count = 46609;
	#10 counter$count = 46610;
	#10 counter$count = 46611;
	#10 counter$count = 46612;
	#10 counter$count = 46613;
	#10 counter$count = 46614;
	#10 counter$count = 46615;
	#10 counter$count = 46616;
	#10 counter$count = 46617;
	#10 counter$count = 46618;
	#10 counter$count = 46619;
	#10 counter$count = 46620;
	#10 counter$count = 46621;
	#10 counter$count = 46622;
	#10 counter$count = 46623;
	#10 counter$count = 46624;
	#10 counter$count = 46625;
	#10 counter$count = 46626;
	#10 counter$count = 46627;
	#10 counter$count = 46628;
	#10 counter$count = 46629;
	#10 counter$count = 46630;
	#10 counter$count = 46631;
	#10 counter$count = 46632;
	#10 counter$count = 46633;
	#10 counter$count = 46634;
	#10 counter$count = 46635;
	#10 counter$count = 46636;
	#10 counter$count = 46637;
	#10 counter$count = 46638;
	#10 counter$count = 46639;
	#10 counter$count = 46640;
	#10 counter$count = 46641;
	#10 counter$count = 46642;
	#10 counter$count = 46643;
	#10 counter$count = 46644;
	#10 counter$count = 46645;
	#10 counter$count = 46646;
	#10 counter$count = 46647;
	#10 counter$count = 46648;
	#10 counter$count = 46649;
	#10 counter$count = 46650;
	#10 counter$count = 46651;
	#10 counter$count = 46652;
	#10 counter$count = 46653;
	#10 counter$count = 46654;
	#10 counter$count = 46655;
	#10 counter$count = 46656;
	#10 counter$count = 46657;
	#10 counter$count = 46658;
	#10 counter$count = 46659;
	#10 counter$count = 46660;
	#10 counter$count = 46661;
	#10 counter$count = 46662;
	#10 counter$count = 46663;
	#10 counter$count = 46664;
	#10 counter$count = 46665;
	#10 counter$count = 46666;
	#10 counter$count = 46667;
	#10 counter$count = 46668;
	#10 counter$count = 46669;
	#10 counter$count = 46670;
	#10 counter$count = 46671;
	#10 counter$count = 46672;
	#10 counter$count = 46673;
	#10 counter$count = 46674;
	#10 counter$count = 46675;
	#10 counter$count = 46676;
	#10 counter$count = 46677;
	#10 counter$count = 46678;
	#10 counter$count = 46679;
	#10 counter$count = 46680;
	#10 counter$count = 46681;
	#10 counter$count = 46682;
	#10 counter$count = 46683;
	#10 counter$count = 46684;
	#10 counter$count = 46685;
	#10 counter$count = 46686;
	#10 counter$count = 46687;
	#10 counter$count = 46688;
	#10 counter$count = 46689;
	#10 counter$count = 46690;
	#10 counter$count = 46691;
	#10 counter$count = 46692;
	#10 counter$count = 46693;
	#10 counter$count = 46694;
	#10 counter$count = 46695;
	#10 counter$count = 46696;
	#10 counter$count = 46697;
	#10 counter$count = 46698;
	#10 counter$count = 46699;
	#10 counter$count = 46700;
	#10 counter$count = 46701;
	#10 counter$count = 46702;
	#10 counter$count = 46703;
	#10 counter$count = 46704;
	#10 counter$count = 46705;
	#10 counter$count = 46706;
	#10 counter$count = 46707;
	#10 counter$count = 46708;
	#10 counter$count = 46709;
	#10 counter$count = 46710;
	#10 counter$count = 46711;
	#10 counter$count = 46712;
	#10 counter$count = 46713;
	#10 counter$count = 46714;
	#10 counter$count = 46715;
	#10 counter$count = 46716;
	#10 counter$count = 46717;
	#10 counter$count = 46718;
	#10 counter$count = 46719;
	#10 counter$count = 46720;
	#10 counter$count = 46721;
	#10 counter$count = 46722;
	#10 counter$count = 46723;
	#10 counter$count = 46724;
	#10 counter$count = 46725;
	#10 counter$count = 46726;
	#10 counter$count = 46727;
	#10 counter$count = 46728;
	#10 counter$count = 46729;
	#10 counter$count = 46730;
	#10 counter$count = 46731;
	#10 counter$count = 46732;
	#10 counter$count = 46733;
	#10 counter$count = 46734;
	#10 counter$count = 46735;
	#10 counter$count = 46736;
	#10 counter$count = 46737;
	#10 counter$count = 46738;
	#10 counter$count = 46739;
	#10 counter$count = 46740;
	#10 counter$count = 46741;
	#10 counter$count = 46742;
	#10 counter$count = 46743;
	#10 counter$count = 46744;
	#10 counter$count = 46745;
	#10 counter$count = 46746;
	#10 counter$count = 46747;
	#10 counter$count = 46748;
	#10 counter$count = 46749;
	#10 counter$count = 46750;
	#10 counter$count = 46751;
	#10 counter$count = 46752;
	#10 counter$count = 46753;
	#10 counter$count = 46754;
	#10 counter$count = 46755;
	#10 counter$count = 46756;
	#10 counter$count = 46757;
	#10 counter$count = 46758;
	#10 counter$count = 46759;
	#10 counter$count = 46760;
	#10 counter$count = 46761;
	#10 counter$count = 46762;
	#10 counter$count = 46763;
	#10 counter$count = 46764;
	#10 counter$count = 46765;
	#10 counter$count = 46766;
	#10 counter$count = 46767;
	#10 counter$count = 46768;
	#10 counter$count = 46769;
	#10 counter$count = 46770;
	#10 counter$count = 46771;
	#10 counter$count = 46772;
	#10 counter$count = 46773;
	#10 counter$count = 46774;
	#10 counter$count = 46775;
	#10 counter$count = 46776;
	#10 counter$count = 46777;
	#10 counter$count = 46778;
	#10 counter$count = 46779;
	#10 counter$count = 46780;
	#10 counter$count = 46781;
	#10 counter$count = 46782;
	#10 counter$count = 46783;
	#10 counter$count = 46784;
	#10 counter$count = 46785;
	#10 counter$count = 46786;
	#10 counter$count = 46787;
	#10 counter$count = 46788;
	#10 counter$count = 46789;
	#10 counter$count = 46790;
	#10 counter$count = 46791;
	#10 counter$count = 46792;
	#10 counter$count = 46793;
	#10 counter$count = 46794;
	#10 counter$count = 46795;
	#10 counter$count = 46796;
	#10 counter$count = 46797;
	#10 counter$count = 46798;
	#10 counter$count = 46799;
	#10 counter$count = 46800;
	#10 counter$count = 46801;
	#10 counter$count = 46802;
	#10 counter$count = 46803;
	#10 counter$count = 46804;
	#10 counter$count = 46805;
	#10 counter$count = 46806;
	#10 counter$count = 46807;
	#10 counter$count = 46808;
	#10 counter$count = 46809;
	#10 counter$count = 46810;
	#10 counter$count = 46811;
	#10 counter$count = 46812;
	#10 counter$count = 46813;
	#10 counter$count = 46814;
	#10 counter$count = 46815;
	#10 counter$count = 46816;
	#10 counter$count = 46817;
	#10 counter$count = 46818;
	#10 counter$count = 46819;
	#10 counter$count = 46820;
	#10 counter$count = 46821;
	#10 counter$count = 46822;
	#10 counter$count = 46823;
	#10 counter$count = 46824;
	#10 counter$count = 46825;
	#10 counter$count = 46826;
	#10 counter$count = 46827;
	#10 counter$count = 46828;
	#10 counter$count = 46829;
	#10 counter$count = 46830;
	#10 counter$count = 46831;
	#10 counter$count = 46832;
	#10 counter$count = 46833;
	#10 counter$count = 46834;
	#10 counter$count = 46835;
	#10 counter$count = 46836;
	#10 counter$count = 46837;
	#10 counter$count = 46838;
	#10 counter$count = 46839;
	#10 counter$count = 46840;
	#10 counter$count = 46841;
	#10 counter$count = 46842;
	#10 counter$count = 46843;
	#10 counter$count = 46844;
	#10 counter$count = 46845;
	#10 counter$count = 46846;
	#10 counter$count = 46847;
	#10 counter$count = 46848;
	#10 counter$count = 46849;
	#10 counter$count = 46850;
	#10 counter$count = 46851;
	#10 counter$count = 46852;
	#10 counter$count = 46853;
	#10 counter$count = 46854;
	#10 counter$count = 46855;
	#10 counter$count = 46856;
	#10 counter$count = 46857;
	#10 counter$count = 46858;
	#10 counter$count = 46859;
	#10 counter$count = 46860;
	#10 counter$count = 46861;
	#10 counter$count = 46862;
	#10 counter$count = 46863;
	#10 counter$count = 46864;
	#10 counter$count = 46865;
	#10 counter$count = 46866;
	#10 counter$count = 46867;
	#10 counter$count = 46868;
	#10 counter$count = 46869;
	#10 counter$count = 46870;
	#10 counter$count = 46871;
	#10 counter$count = 46872;
	#10 counter$count = 46873;
	#10 counter$count = 46874;
	#10 counter$count = 46875;
	#10 counter$count = 46876;
	#10 counter$count = 46877;
	#10 counter$count = 46878;
	#10 counter$count = 46879;
	#10 counter$count = 46880;
	#10 counter$count = 46881;
	#10 counter$count = 46882;
	#10 counter$count = 46883;
	#10 counter$count = 46884;
	#10 counter$count = 46885;
	#10 counter$count = 46886;
	#10 counter$count = 46887;
	#10 counter$count = 46888;
	#10 counter$count = 46889;
	#10 counter$count = 46890;
	#10 counter$count = 46891;
	#10 counter$count = 46892;
	#10 counter$count = 46893;
	#10 counter$count = 46894;
	#10 counter$count = 46895;
	#10 counter$count = 46896;
	#10 counter$count = 46897;
	#10 counter$count = 46898;
	#10 counter$count = 46899;
	#10 counter$count = 46900;
	#10 counter$count = 46901;
	#10 counter$count = 46902;
	#10 counter$count = 46903;
	#10 counter$count = 46904;
	#10 counter$count = 46905;
	#10 counter$count = 46906;
	#10 counter$count = 46907;
	#10 counter$count = 46908;
	#10 counter$count = 46909;
	#10 counter$count = 46910;
	#10 counter$count = 46911;
	#10 counter$count = 46912;
	#10 counter$count = 46913;
	#10 counter$count = 46914;
	#10 counter$count = 46915;
	#10 counter$count = 46916;
	#10 counter$count = 46917;
	#10 counter$count = 46918;
	#10 counter$count = 46919;
	#10 counter$count = 46920;
	#10 counter$count = 46921;
	#10 counter$count = 46922;
	#10 counter$count = 46923;
	#10 counter$count = 46924;
	#10 counter$count = 46925;
	#10 counter$count = 46926;
	#10 counter$count = 46927;
	#10 counter$count = 46928;
	#10 counter$count = 46929;
	#10 counter$count = 46930;
	#10 counter$count = 46931;
	#10 counter$count = 46932;
	#10 counter$count = 46933;
	#10 counter$count = 46934;
	#10 counter$count = 46935;
	#10 counter$count = 46936;
	#10 counter$count = 46937;
	#10 counter$count = 46938;
	#10 counter$count = 46939;
	#10 counter$count = 46940;
	#10 counter$count = 46941;
	#10 counter$count = 46942;
	#10 counter$count = 46943;
	#10 counter$count = 46944;
	#10 counter$count = 46945;
	#10 counter$count = 46946;
	#10 counter$count = 46947;
	#10 counter$count = 46948;
	#10 counter$count = 46949;
	#10 counter$count = 46950;
	#10 counter$count = 46951;
	#10 counter$count = 46952;
	#10 counter$count = 46953;
	#10 counter$count = 46954;
	#10 counter$count = 46955;
	#10 counter$count = 46956;
	#10 counter$count = 46957;
	#10 counter$count = 46958;
	#10 counter$count = 46959;
	#10 counter$count = 46960;
	#10 counter$count = 46961;
	#10 counter$count = 46962;
	#10 counter$count = 46963;
	#10 counter$count = 46964;
	#10 counter$count = 46965;
	#10 counter$count = 46966;
	#10 counter$count = 46967;
	#10 counter$count = 46968;
	#10 counter$count = 46969;
	#10 counter$count = 46970;
	#10 counter$count = 46971;
	#10 counter$count = 46972;
	#10 counter$count = 46973;
	#10 counter$count = 46974;
	#10 counter$count = 46975;
	#10 counter$count = 46976;
	#10 counter$count = 46977;
	#10 counter$count = 46978;
	#10 counter$count = 46979;
	#10 counter$count = 46980;
	#10 counter$count = 46981;
	#10 counter$count = 46982;
	#10 counter$count = 46983;
	#10 counter$count = 46984;
	#10 counter$count = 46985;
	#10 counter$count = 46986;
	#10 counter$count = 46987;
	#10 counter$count = 46988;
	#10 counter$count = 46989;
	#10 counter$count = 46990;
	#10 counter$count = 46991;
	#10 counter$count = 46992;
	#10 counter$count = 46993;
	#10 counter$count = 46994;
	#10 counter$count = 46995;
	#10 counter$count = 46996;
	#10 counter$count = 46997;
	#10 counter$count = 46998;
	#10 counter$count = 46999;
	#10 counter$count = 47000;
	#10 counter$count = 47001;
	#10 counter$count = 47002;
	#10 counter$count = 47003;
	#10 counter$count = 47004;
	#10 counter$count = 47005;
	#10 counter$count = 47006;
	#10 counter$count = 47007;
	#10 counter$count = 47008;
	#10 counter$count = 47009;
	#10 counter$count = 47010;
	#10 counter$count = 47011;
	#10 counter$count = 47012;
	#10 counter$count = 47013;
	#10 counter$count = 47014;
	#10 counter$count = 47015;
	#10 counter$count = 47016;
	#10 counter$count = 47017;
	#10 counter$count = 47018;
	#10 counter$count = 47019;
	#10 counter$count = 47020;
	#10 counter$count = 47021;
	#10 counter$count = 47022;
	#10 counter$count = 47023;
	#10 counter$count = 47024;
	#10 counter$count = 47025;
	#10 counter$count = 47026;
	#10 counter$count = 47027;
	#10 counter$count = 47028;
	#10 counter$count = 47029;
	#10 counter$count = 47030;
	#10 counter$count = 47031;
	#10 counter$count = 47032;
	#10 counter$count = 47033;
	#10 counter$count = 47034;
	#10 counter$count = 47035;
	#10 counter$count = 47036;
	#10 counter$count = 47037;
	#10 counter$count = 47038;
	#10 counter$count = 47039;
	#10 counter$count = 47040;
	#10 counter$count = 47041;
	#10 counter$count = 47042;
	#10 counter$count = 47043;
	#10 counter$count = 47044;
	#10 counter$count = 47045;
	#10 counter$count = 47046;
	#10 counter$count = 47047;
	#10 counter$count = 47048;
	#10 counter$count = 47049;
	#10 counter$count = 47050;
	#10 counter$count = 47051;
	#10 counter$count = 47052;
	#10 counter$count = 47053;
	#10 counter$count = 47054;
	#10 counter$count = 47055;
	#10 counter$count = 47056;
	#10 counter$count = 47057;
	#10 counter$count = 47058;
	#10 counter$count = 47059;
	#10 counter$count = 47060;
	#10 counter$count = 47061;
	#10 counter$count = 47062;
	#10 counter$count = 47063;
	#10 counter$count = 47064;
	#10 counter$count = 47065;
	#10 counter$count = 47066;
	#10 counter$count = 47067;
	#10 counter$count = 47068;
	#10 counter$count = 47069;
	#10 counter$count = 47070;
	#10 counter$count = 47071;
	#10 counter$count = 47072;
	#10 counter$count = 47073;
	#10 counter$count = 47074;
	#10 counter$count = 47075;
	#10 counter$count = 47076;
	#10 counter$count = 47077;
	#10 counter$count = 47078;
	#10 counter$count = 47079;
	#10 counter$count = 47080;
	#10 counter$count = 47081;
	#10 counter$count = 47082;
	#10 counter$count = 47083;
	#10 counter$count = 47084;
	#10 counter$count = 47085;
	#10 counter$count = 47086;
	#10 counter$count = 47087;
	#10 counter$count = 47088;
	#10 counter$count = 47089;
	#10 counter$count = 47090;
	#10 counter$count = 47091;
	#10 counter$count = 47092;
	#10 counter$count = 47093;
	#10 counter$count = 47094;
	#10 counter$count = 47095;
	#10 counter$count = 47096;
	#10 counter$count = 47097;
	#10 counter$count = 47098;
	#10 counter$count = 47099;
	#10 counter$count = 47100;
	#10 counter$count = 47101;
	#10 counter$count = 47102;
	#10 counter$count = 47103;
	#10 counter$count = 47104;
	#10 counter$count = 47105;
	#10 counter$count = 47106;
	#10 counter$count = 47107;
	#10 counter$count = 47108;
	#10 counter$count = 47109;
	#10 counter$count = 47110;
	#10 counter$count = 47111;
	#10 counter$count = 47112;
	#10 counter$count = 47113;
	#10 counter$count = 47114;
	#10 counter$count = 47115;
	#10 counter$count = 47116;
	#10 counter$count = 47117;
	#10 counter$count = 47118;
	#10 counter$count = 47119;
	#10 counter$count = 47120;
	#10 counter$count = 47121;
	#10 counter$count = 47122;
	#10 counter$count = 47123;
	#10 counter$count = 47124;
	#10 counter$count = 47125;
	#10 counter$count = 47126;
	#10 counter$count = 47127;
	#10 counter$count = 47128;
	#10 counter$count = 47129;
	#10 counter$count = 47130;
	#10 counter$count = 47131;
	#10 counter$count = 47132;
	#10 counter$count = 47133;
	#10 counter$count = 47134;
	#10 counter$count = 47135;
	#10 counter$count = 47136;
	#10 counter$count = 47137;
	#10 counter$count = 47138;
	#10 counter$count = 47139;
	#10 counter$count = 47140;
	#10 counter$count = 47141;
	#10 counter$count = 47142;
	#10 counter$count = 47143;
	#10 counter$count = 47144;
	#10 counter$count = 47145;
	#10 counter$count = 47146;
	#10 counter$count = 47147;
	#10 counter$count = 47148;
	#10 counter$count = 47149;
	#10 counter$count = 47150;
	#10 counter$count = 47151;
	#10 counter$count = 47152;
	#10 counter$count = 47153;
	#10 counter$count = 47154;
	#10 counter$count = 47155;
	#10 counter$count = 47156;
	#10 counter$count = 47157;
	#10 counter$count = 47158;
	#10 counter$count = 47159;
	#10 counter$count = 47160;
	#10 counter$count = 47161;
	#10 counter$count = 47162;
	#10 counter$count = 47163;
	#10 counter$count = 47164;
	#10 counter$count = 47165;
	#10 counter$count = 47166;
	#10 counter$count = 47167;
	#10 counter$count = 47168;
	#10 counter$count = 47169;
	#10 counter$count = 47170;
	#10 counter$count = 47171;
	#10 counter$count = 47172;
	#10 counter$count = 47173;
	#10 counter$count = 47174;
	#10 counter$count = 47175;
	#10 counter$count = 47176;
	#10 counter$count = 47177;
	#10 counter$count = 47178;
	#10 counter$count = 47179;
	#10 counter$count = 47180;
	#10 counter$count = 47181;
	#10 counter$count = 47182;
	#10 counter$count = 47183;
	#10 counter$count = 47184;
	#10 counter$count = 47185;
	#10 counter$count = 47186;
	#10 counter$count = 47187;
	#10 counter$count = 47188;
	#10 counter$count = 47189;
	#10 counter$count = 47190;
	#10 counter$count = 47191;
	#10 counter$count = 47192;
	#10 counter$count = 47193;
	#10 counter$count = 47194;
	#10 counter$count = 47195;
	#10 counter$count = 47196;
	#10 counter$count = 47197;
	#10 counter$count = 47198;
	#10 counter$count = 47199;
	#10 counter$count = 47200;
	#10 counter$count = 47201;
	#10 counter$count = 47202;
	#10 counter$count = 47203;
	#10 counter$count = 47204;
	#10 counter$count = 47205;
	#10 counter$count = 47206;
	#10 counter$count = 47207;
	#10 counter$count = 47208;
	#10 counter$count = 47209;
	#10 counter$count = 47210;
	#10 counter$count = 47211;
	#10 counter$count = 47212;
	#10 counter$count = 47213;
	#10 counter$count = 47214;
	#10 counter$count = 47215;
	#10 counter$count = 47216;
	#10 counter$count = 47217;
	#10 counter$count = 47218;
	#10 counter$count = 47219;
	#10 counter$count = 47220;
	#10 counter$count = 47221;
	#10 counter$count = 47222;
	#10 counter$count = 47223;
	#10 counter$count = 47224;
	#10 counter$count = 47225;
	#10 counter$count = 47226;
	#10 counter$count = 47227;
	#10 counter$count = 47228;
	#10 counter$count = 47229;
	#10 counter$count = 47230;
	#10 counter$count = 47231;
	#10 counter$count = 47232;
	#10 counter$count = 47233;
	#10 counter$count = 47234;
	#10 counter$count = 47235;
	#10 counter$count = 47236;
	#10 counter$count = 47237;
	#10 counter$count = 47238;
	#10 counter$count = 47239;
	#10 counter$count = 47240;
	#10 counter$count = 47241;
	#10 counter$count = 47242;
	#10 counter$count = 47243;
	#10 counter$count = 47244;
	#10 counter$count = 47245;
	#10 counter$count = 47246;
	#10 counter$count = 47247;
	#10 counter$count = 47248;
	#10 counter$count = 47249;
	#10 counter$count = 47250;
	#10 counter$count = 47251;
	#10 counter$count = 47252;
	#10 counter$count = 47253;
	#10 counter$count = 47254;
	#10 counter$count = 47255;
	#10 counter$count = 47256;
	#10 counter$count = 47257;
	#10 counter$count = 47258;
	#10 counter$count = 47259;
	#10 counter$count = 47260;
	#10 counter$count = 47261;
	#10 counter$count = 47262;
	#10 counter$count = 47263;
	#10 counter$count = 47264;
	#10 counter$count = 47265;
	#10 counter$count = 47266;
	#10 counter$count = 47267;
	#10 counter$count = 47268;
	#10 counter$count = 47269;
	#10 counter$count = 47270;
	#10 counter$count = 47271;
	#10 counter$count = 47272;
	#10 counter$count = 47273;
	#10 counter$count = 47274;
	#10 counter$count = 47275;
	#10 counter$count = 47276;
	#10 counter$count = 47277;
	#10 counter$count = 47278;
	#10 counter$count = 47279;
	#10 counter$count = 47280;
	#10 counter$count = 47281;
	#10 counter$count = 47282;
	#10 counter$count = 47283;
	#10 counter$count = 47284;
	#10 counter$count = 47285;
	#10 counter$count = 47286;
	#10 counter$count = 47287;
	#10 counter$count = 47288;
	#10 counter$count = 47289;
	#10 counter$count = 47290;
	#10 counter$count = 47291;
	#10 counter$count = 47292;
	#10 counter$count = 47293;
	#10 counter$count = 47294;
	#10 counter$count = 47295;
	#10 counter$count = 47296;
	#10 counter$count = 47297;
	#10 counter$count = 47298;
	#10 counter$count = 47299;
	#10 counter$count = 47300;
	#10 counter$count = 47301;
	#10 counter$count = 47302;
	#10 counter$count = 47303;
	#10 counter$count = 47304;
	#10 counter$count = 47305;
	#10 counter$count = 47306;
	#10 counter$count = 47307;
	#10 counter$count = 47308;
	#10 counter$count = 47309;
	#10 counter$count = 47310;
	#10 counter$count = 47311;
	#10 counter$count = 47312;
	#10 counter$count = 47313;
	#10 counter$count = 47314;
	#10 counter$count = 47315;
	#10 counter$count = 47316;
	#10 counter$count = 47317;
	#10 counter$count = 47318;
	#10 counter$count = 47319;
	#10 counter$count = 47320;
	#10 counter$count = 47321;
	#10 counter$count = 47322;
	#10 counter$count = 47323;
	#10 counter$count = 47324;
	#10 counter$count = 47325;
	#10 counter$count = 47326;
	#10 counter$count = 47327;
	#10 counter$count = 47328;
	#10 counter$count = 47329;
	#10 counter$count = 47330;
	#10 counter$count = 47331;
	#10 counter$count = 47332;
	#10 counter$count = 47333;
	#10 counter$count = 47334;
	#10 counter$count = 47335;
	#10 counter$count = 47336;
	#10 counter$count = 47337;
	#10 counter$count = 47338;
	#10 counter$count = 47339;
	#10 counter$count = 47340;
	#10 counter$count = 47341;
	#10 counter$count = 47342;
	#10 counter$count = 47343;
	#10 counter$count = 47344;
	#10 counter$count = 47345;
	#10 counter$count = 47346;
	#10 counter$count = 47347;
	#10 counter$count = 47348;
	#10 counter$count = 47349;
	#10 counter$count = 47350;
	#10 counter$count = 47351;
	#10 counter$count = 47352;
	#10 counter$count = 47353;
	#10 counter$count = 47354;
	#10 counter$count = 47355;
	#10 counter$count = 47356;
	#10 counter$count = 47357;
	#10 counter$count = 47358;
	#10 counter$count = 47359;
	#10 counter$count = 47360;
	#10 counter$count = 47361;
	#10 counter$count = 47362;
	#10 counter$count = 47363;
	#10 counter$count = 47364;
	#10 counter$count = 47365;
	#10 counter$count = 47366;
	#10 counter$count = 47367;
	#10 counter$count = 47368;
	#10 counter$count = 47369;
	#10 counter$count = 47370;
	#10 counter$count = 47371;
	#10 counter$count = 47372;
	#10 counter$count = 47373;
	#10 counter$count = 47374;
	#10 counter$count = 47375;
	#10 counter$count = 47376;
	#10 counter$count = 47377;
	#10 counter$count = 47378;
	#10 counter$count = 47379;
	#10 counter$count = 47380;
	#10 counter$count = 47381;
	#10 counter$count = 47382;
	#10 counter$count = 47383;
	#10 counter$count = 47384;
	#10 counter$count = 47385;
	#10 counter$count = 47386;
	#10 counter$count = 47387;
	#10 counter$count = 47388;
	#10 counter$count = 47389;
	#10 counter$count = 47390;
	#10 counter$count = 47391;
	#10 counter$count = 47392;
	#10 counter$count = 47393;
	#10 counter$count = 47394;
	#10 counter$count = 47395;
	#10 counter$count = 47396;
	#10 counter$count = 47397;
	#10 counter$count = 47398;
	#10 counter$count = 47399;
	#10 counter$count = 47400;
	#10 counter$count = 47401;
	#10 counter$count = 47402;
	#10 counter$count = 47403;
	#10 counter$count = 47404;
	#10 counter$count = 47405;
	#10 counter$count = 47406;
	#10 counter$count = 47407;
	#10 counter$count = 47408;
	#10 counter$count = 47409;
	#10 counter$count = 47410;
	#10 counter$count = 47411;
	#10 counter$count = 47412;
	#10 counter$count = 47413;
	#10 counter$count = 47414;
	#10 counter$count = 47415;
	#10 counter$count = 47416;
	#10 counter$count = 47417;
	#10 counter$count = 47418;
	#10 counter$count = 47419;
	#10 counter$count = 47420;
	#10 counter$count = 47421;
	#10 counter$count = 47422;
	#10 counter$count = 47423;
	#10 counter$count = 47424;
	#10 counter$count = 47425;
	#10 counter$count = 47426;
	#10 counter$count = 47427;
	#10 counter$count = 47428;
	#10 counter$count = 47429;
	#10 counter$count = 47430;
	#10 counter$count = 47431;
	#10 counter$count = 47432;
	#10 counter$count = 47433;
	#10 counter$count = 47434;
	#10 counter$count = 47435;
	#10 counter$count = 47436;
	#10 counter$count = 47437;
	#10 counter$count = 47438;
	#10 counter$count = 47439;
	#10 counter$count = 47440;
	#10 counter$count = 47441;
	#10 counter$count = 47442;
	#10 counter$count = 47443;
	#10 counter$count = 47444;
	#10 counter$count = 47445;
	#10 counter$count = 47446;
	#10 counter$count = 47447;
	#10 counter$count = 47448;
	#10 counter$count = 47449;
	#10 counter$count = 47450;
	#10 counter$count = 47451;
	#10 counter$count = 47452;
	#10 counter$count = 47453;
	#10 counter$count = 47454;
	#10 counter$count = 47455;
	#10 counter$count = 47456;
	#10 counter$count = 47457;
	#10 counter$count = 47458;
	#10 counter$count = 47459;
	#10 counter$count = 47460;
	#10 counter$count = 47461;
	#10 counter$count = 47462;
	#10 counter$count = 47463;
	#10 counter$count = 47464;
	#10 counter$count = 47465;
	#10 counter$count = 47466;
	#10 counter$count = 47467;
	#10 counter$count = 47468;
	#10 counter$count = 47469;
	#10 counter$count = 47470;
	#10 counter$count = 47471;
	#10 counter$count = 47472;
	#10 counter$count = 47473;
	#10 counter$count = 47474;
	#10 counter$count = 47475;
	#10 counter$count = 47476;
	#10 counter$count = 47477;
	#10 counter$count = 47478;
	#10 counter$count = 47479;
	#10 counter$count = 47480;
	#10 counter$count = 47481;
	#10 counter$count = 47482;
	#10 counter$count = 47483;
	#10 counter$count = 47484;
	#10 counter$count = 47485;
	#10 counter$count = 47486;
	#10 counter$count = 47487;
	#10 counter$count = 47488;
	#10 counter$count = 47489;
	#10 counter$count = 47490;
	#10 counter$count = 47491;
	#10 counter$count = 47492;
	#10 counter$count = 47493;
	#10 counter$count = 47494;
	#10 counter$count = 47495;
	#10 counter$count = 47496;
	#10 counter$count = 47497;
	#10 counter$count = 47498;
	#10 counter$count = 47499;
	#10 counter$count = 47500;
	#10 counter$count = 47501;
	#10 counter$count = 47502;
	#10 counter$count = 47503;
	#10 counter$count = 47504;
	#10 counter$count = 47505;
	#10 counter$count = 47506;
	#10 counter$count = 47507;
	#10 counter$count = 47508;
	#10 counter$count = 47509;
	#10 counter$count = 47510;
	#10 counter$count = 47511;
	#10 counter$count = 47512;
	#10 counter$count = 47513;
	#10 counter$count = 47514;
	#10 counter$count = 47515;
	#10 counter$count = 47516;
	#10 counter$count = 47517;
	#10 counter$count = 47518;
	#10 counter$count = 47519;
	#10 counter$count = 47520;
	#10 counter$count = 47521;
	#10 counter$count = 47522;
	#10 counter$count = 47523;
	#10 counter$count = 47524;
	#10 counter$count = 47525;
	#10 counter$count = 47526;
	#10 counter$count = 47527;
	#10 counter$count = 47528;
	#10 counter$count = 47529;
	#10 counter$count = 47530;
	#10 counter$count = 47531;
	#10 counter$count = 47532;
	#10 counter$count = 47533;
	#10 counter$count = 47534;
	#10 counter$count = 47535;
	#10 counter$count = 47536;
	#10 counter$count = 47537;
	#10 counter$count = 47538;
	#10 counter$count = 47539;
	#10 counter$count = 47540;
	#10 counter$count = 47541;
	#10 counter$count = 47542;
	#10 counter$count = 47543;
	#10 counter$count = 47544;
	#10 counter$count = 47545;
	#10 counter$count = 47546;
	#10 counter$count = 47547;
	#10 counter$count = 47548;
	#10 counter$count = 47549;
	#10 counter$count = 47550;
	#10 counter$count = 47551;
	#10 counter$count = 47552;
	#10 counter$count = 47553;
	#10 counter$count = 47554;
	#10 counter$count = 47555;
	#10 counter$count = 47556;
	#10 counter$count = 47557;
	#10 counter$count = 47558;
	#10 counter$count = 47559;
	#10 counter$count = 47560;
	#10 counter$count = 47561;
	#10 counter$count = 47562;
	#10 counter$count = 47563;
	#10 counter$count = 47564;
	#10 counter$count = 47565;
	#10 counter$count = 47566;
	#10 counter$count = 47567;
	#10 counter$count = 47568;
	#10 counter$count = 47569;
	#10 counter$count = 47570;
	#10 counter$count = 47571;
	#10 counter$count = 47572;
	#10 counter$count = 47573;
	#10 counter$count = 47574;
	#10 counter$count = 47575;
	#10 counter$count = 47576;
	#10 counter$count = 47577;
	#10 counter$count = 47578;
	#10 counter$count = 47579;
	#10 counter$count = 47580;
	#10 counter$count = 47581;
	#10 counter$count = 47582;
	#10 counter$count = 47583;
	#10 counter$count = 47584;
	#10 counter$count = 47585;
	#10 counter$count = 47586;
	#10 counter$count = 47587;
	#10 counter$count = 47588;
	#10 counter$count = 47589;
	#10 counter$count = 47590;
	#10 counter$count = 47591;
	#10 counter$count = 47592;
	#10 counter$count = 47593;
	#10 counter$count = 47594;
	#10 counter$count = 47595;
	#10 counter$count = 47596;
	#10 counter$count = 47597;
	#10 counter$count = 47598;
	#10 counter$count = 47599;
	#10 counter$count = 47600;
	#10 counter$count = 47601;
	#10 counter$count = 47602;
	#10 counter$count = 47603;
	#10 counter$count = 47604;
	#10 counter$count = 47605;
	#10 counter$count = 47606;
	#10 counter$count = 47607;
	#10 counter$count = 47608;
	#10 counter$count = 47609;
	#10 counter$count = 47610;
	#10 counter$count = 47611;
	#10 counter$count = 47612;
	#10 counter$count = 47613;
	#10 counter$count = 47614;
	#10 counter$count = 47615;
	#10 counter$count = 47616;
	#10 counter$count = 47617;
	#10 counter$count = 47618;
	#10 counter$count = 47619;
	#10 counter$count = 47620;
	#10 counter$count = 47621;
	#10 counter$count = 47622;
	#10 counter$count = 47623;
	#10 counter$count = 47624;
	#10 counter$count = 47625;
	#10 counter$count = 47626;
	#10 counter$count = 47627;
	#10 counter$count = 47628;
	#10 counter$count = 47629;
	#10 counter$count = 47630;
	#10 counter$count = 47631;
	#10 counter$count = 47632;
	#10 counter$count = 47633;
	#10 counter$count = 47634;
	#10 counter$count = 47635;
	#10 counter$count = 47636;
	#10 counter$count = 47637;
	#10 counter$count = 47638;
	#10 counter$count = 47639;
	#10 counter$count = 47640;
	#10 counter$count = 47641;
	#10 counter$count = 47642;
	#10 counter$count = 47643;
	#10 counter$count = 47644;
	#10 counter$count = 47645;
	#10 counter$count = 47646;
	#10 counter$count = 47647;
	#10 counter$count = 47648;
	#10 counter$count = 47649;
	#10 counter$count = 47650;
	#10 counter$count = 47651;
	#10 counter$count = 47652;
	#10 counter$count = 47653;
	#10 counter$count = 47654;
	#10 counter$count = 47655;
	#10 counter$count = 47656;
	#10 counter$count = 47657;
	#10 counter$count = 47658;
	#10 counter$count = 47659;
	#10 counter$count = 47660;
	#10 counter$count = 47661;
	#10 counter$count = 47662;
	#10 counter$count = 47663;
	#10 counter$count = 47664;
	#10 counter$count = 47665;
	#10 counter$count = 47666;
	#10 counter$count = 47667;
	#10 counter$count = 47668;
	#10 counter$count = 47669;
	#10 counter$count = 47670;
	#10 counter$count = 47671;
	#10 counter$count = 47672;
	#10 counter$count = 47673;
	#10 counter$count = 47674;
	#10 counter$count = 47675;
	#10 counter$count = 47676;
	#10 counter$count = 47677;
	#10 counter$count = 47678;
	#10 counter$count = 47679;
	#10 counter$count = 47680;
	#10 counter$count = 47681;
	#10 counter$count = 47682;
	#10 counter$count = 47683;
	#10 counter$count = 47684;
	#10 counter$count = 47685;
	#10 counter$count = 47686;
	#10 counter$count = 47687;
	#10 counter$count = 47688;
	#10 counter$count = 47689;
	#10 counter$count = 47690;
	#10 counter$count = 47691;
	#10 counter$count = 47692;
	#10 counter$count = 47693;
	#10 counter$count = 47694;
	#10 counter$count = 47695;
	#10 counter$count = 47696;
	#10 counter$count = 47697;
	#10 counter$count = 47698;
	#10 counter$count = 47699;
	#10 counter$count = 47700;
	#10 counter$count = 47701;
	#10 counter$count = 47702;
	#10 counter$count = 47703;
	#10 counter$count = 47704;
	#10 counter$count = 47705;
	#10 counter$count = 47706;
	#10 counter$count = 47707;
	#10 counter$count = 47708;
	#10 counter$count = 47709;
	#10 counter$count = 47710;
	#10 counter$count = 47711;
	#10 counter$count = 47712;
	#10 counter$count = 47713;
	#10 counter$count = 47714;
	#10 counter$count = 47715;
	#10 counter$count = 47716;
	#10 counter$count = 47717;
	#10 counter$count = 47718;
	#10 counter$count = 47719;
	#10 counter$count = 47720;
	#10 counter$count = 47721;
	#10 counter$count = 47722;
	#10 counter$count = 47723;
	#10 counter$count = 47724;
	#10 counter$count = 47725;
	#10 counter$count = 47726;
	#10 counter$count = 47727;
	#10 counter$count = 47728;
	#10 counter$count = 47729;
	#10 counter$count = 47730;
	#10 counter$count = 47731;
	#10 counter$count = 47732;
	#10 counter$count = 47733;
	#10 counter$count = 47734;
	#10 counter$count = 47735;
	#10 counter$count = 47736;
	#10 counter$count = 47737;
	#10 counter$count = 47738;
	#10 counter$count = 47739;
	#10 counter$count = 47740;
	#10 counter$count = 47741;
	#10 counter$count = 47742;
	#10 counter$count = 47743;
	#10 counter$count = 47744;
	#10 counter$count = 47745;
	#10 counter$count = 47746;
	#10 counter$count = 47747;
	#10 counter$count = 47748;
	#10 counter$count = 47749;
	#10 counter$count = 47750;
	#10 counter$count = 47751;
	#10 counter$count = 47752;
	#10 counter$count = 47753;
	#10 counter$count = 47754;
	#10 counter$count = 47755;
	#10 counter$count = 47756;
	#10 counter$count = 47757;
	#10 counter$count = 47758;
	#10 counter$count = 47759;
	#10 counter$count = 47760;
	#10 counter$count = 47761;
	#10 counter$count = 47762;
	#10 counter$count = 47763;
	#10 counter$count = 47764;
	#10 counter$count = 47765;
	#10 counter$count = 47766;
	#10 counter$count = 47767;
	#10 counter$count = 47768;
	#10 counter$count = 47769;
	#10 counter$count = 47770;
	#10 counter$count = 47771;
	#10 counter$count = 47772;
	#10 counter$count = 47773;
	#10 counter$count = 47774;
	#10 counter$count = 47775;
	#10 counter$count = 47776;
	#10 counter$count = 47777;
	#10 counter$count = 47778;
	#10 counter$count = 47779;
	#10 counter$count = 47780;
	#10 counter$count = 47781;
	#10 counter$count = 47782;
	#10 counter$count = 47783;
	#10 counter$count = 47784;
	#10 counter$count = 47785;
	#10 counter$count = 47786;
	#10 counter$count = 47787;
	#10 counter$count = 47788;
	#10 counter$count = 47789;
	#10 counter$count = 47790;
	#10 counter$count = 47791;
	#10 counter$count = 47792;
	#10 counter$count = 47793;
	#10 counter$count = 47794;
	#10 counter$count = 47795;
	#10 counter$count = 47796;
	#10 counter$count = 47797;
	#10 counter$count = 47798;
	#10 counter$count = 47799;
	#10 counter$count = 47800;
	#10 counter$count = 47801;
	#10 counter$count = 47802;
	#10 counter$count = 47803;
	#10 counter$count = 47804;
	#10 counter$count = 47805;
	#10 counter$count = 47806;
	#10 counter$count = 47807;
	#10 counter$count = 47808;
	#10 counter$count = 47809;
	#10 counter$count = 47810;
	#10 counter$count = 47811;
	#10 counter$count = 47812;
	#10 counter$count = 47813;
	#10 counter$count = 47814;
	#10 counter$count = 47815;
	#10 counter$count = 47816;
	#10 counter$count = 47817;
	#10 counter$count = 47818;
	#10 counter$count = 47819;
	#10 counter$count = 47820;
	#10 counter$count = 47821;
	#10 counter$count = 47822;
	#10 counter$count = 47823;
	#10 counter$count = 47824;
	#10 counter$count = 47825;
	#10 counter$count = 47826;
	#10 counter$count = 47827;
	#10 counter$count = 47828;
	#10 counter$count = 47829;
	#10 counter$count = 47830;
	#10 counter$count = 47831;
	#10 counter$count = 47832;
	#10 counter$count = 47833;
	#10 counter$count = 47834;
	#10 counter$count = 47835;
	#10 counter$count = 47836;
	#10 counter$count = 47837;
	#10 counter$count = 47838;
	#10 counter$count = 47839;
	#10 counter$count = 47840;
	#10 counter$count = 47841;
	#10 counter$count = 47842;
	#10 counter$count = 47843;
	#10 counter$count = 47844;
	#10 counter$count = 47845;
	#10 counter$count = 47846;
	#10 counter$count = 47847;
	#10 counter$count = 47848;
	#10 counter$count = 47849;
	#10 counter$count = 47850;
	#10 counter$count = 47851;
	#10 counter$count = 47852;
	#10 counter$count = 47853;
	#10 counter$count = 47854;
	#10 counter$count = 47855;
	#10 counter$count = 47856;
	#10 counter$count = 47857;
	#10 counter$count = 47858;
	#10 counter$count = 47859;
	#10 counter$count = 47860;
	#10 counter$count = 47861;
	#10 counter$count = 47862;
	#10 counter$count = 47863;
	#10 counter$count = 47864;
	#10 counter$count = 47865;
	#10 counter$count = 47866;
	#10 counter$count = 47867;
	#10 counter$count = 47868;
	#10 counter$count = 47869;
	#10 counter$count = 47870;
	#10 counter$count = 47871;
	#10 counter$count = 47872;
	#10 counter$count = 47873;
	#10 counter$count = 47874;
	#10 counter$count = 47875;
	#10 counter$count = 47876;
	#10 counter$count = 47877;
	#10 counter$count = 47878;
	#10 counter$count = 47879;
	#10 counter$count = 47880;
	#10 counter$count = 47881;
	#10 counter$count = 47882;
	#10 counter$count = 47883;
	#10 counter$count = 47884;
	#10 counter$count = 47885;
	#10 counter$count = 47886;
	#10 counter$count = 47887;
	#10 counter$count = 47888;
	#10 counter$count = 47889;
	#10 counter$count = 47890;
	#10 counter$count = 47891;
	#10 counter$count = 47892;
	#10 counter$count = 47893;
	#10 counter$count = 47894;
	#10 counter$count = 47895;
	#10 counter$count = 47896;
	#10 counter$count = 47897;
	#10 counter$count = 47898;
	#10 counter$count = 47899;
	#10 counter$count = 47900;
	#10 counter$count = 47901;
	#10 counter$count = 47902;
	#10 counter$count = 47903;
	#10 counter$count = 47904;
	#10 counter$count = 47905;
	#10 counter$count = 47906;
	#10 counter$count = 47907;
	#10 counter$count = 47908;
	#10 counter$count = 47909;
	#10 counter$count = 47910;
	#10 counter$count = 47911;
	#10 counter$count = 47912;
	#10 counter$count = 47913;
	#10 counter$count = 47914;
	#10 counter$count = 47915;
	#10 counter$count = 47916;
	#10 counter$count = 47917;
	#10 counter$count = 47918;
	#10 counter$count = 47919;
	#10 counter$count = 47920;
	#10 counter$count = 47921;
	#10 counter$count = 47922;
	#10 counter$count = 47923;
	#10 counter$count = 47924;
	#10 counter$count = 47925;
	#10 counter$count = 47926;
	#10 counter$count = 47927;
	#10 counter$count = 47928;
	#10 counter$count = 47929;
	#10 counter$count = 47930;
	#10 counter$count = 47931;
	#10 counter$count = 47932;
	#10 counter$count = 47933;
	#10 counter$count = 47934;
	#10 counter$count = 47935;
	#10 counter$count = 47936;
	#10 counter$count = 47937;
	#10 counter$count = 47938;
	#10 counter$count = 47939;
	#10 counter$count = 47940;
	#10 counter$count = 47941;
	#10 counter$count = 47942;
	#10 counter$count = 47943;
	#10 counter$count = 47944;
	#10 counter$count = 47945;
	#10 counter$count = 47946;
	#10 counter$count = 47947;
	#10 counter$count = 47948;
	#10 counter$count = 47949;
	#10 counter$count = 47950;
	#10 counter$count = 47951;
	#10 counter$count = 47952;
	#10 counter$count = 47953;
	#10 counter$count = 47954;
	#10 counter$count = 47955;
	#10 counter$count = 47956;
	#10 counter$count = 47957;
	#10 counter$count = 47958;
	#10 counter$count = 47959;
	#10 counter$count = 47960;
	#10 counter$count = 47961;
	#10 counter$count = 47962;
	#10 counter$count = 47963;
	#10 counter$count = 47964;
	#10 counter$count = 47965;
	#10 counter$count = 47966;
	#10 counter$count = 47967;
	#10 counter$count = 47968;
	#10 counter$count = 47969;
	#10 counter$count = 47970;
	#10 counter$count = 47971;
	#10 counter$count = 47972;
	#10 counter$count = 47973;
	#10 counter$count = 47974;
	#10 counter$count = 47975;
	#10 counter$count = 47976;
	#10 counter$count = 47977;
	#10 counter$count = 47978;
	#10 counter$count = 47979;
	#10 counter$count = 47980;
	#10 counter$count = 47981;
	#10 counter$count = 47982;
	#10 counter$count = 47983;
	#10 counter$count = 47984;
	#10 counter$count = 47985;
	#10 counter$count = 47986;
	#10 counter$count = 47987;
	#10 counter$count = 47988;
	#10 counter$count = 47989;
	#10 counter$count = 47990;
	#10 counter$count = 47991;
	#10 counter$count = 47992;
	#10 counter$count = 47993;
	#10 counter$count = 47994;
	#10 counter$count = 47995;
	#10 counter$count = 47996;
	#10 counter$count = 47997;
	#10 counter$count = 47998;
	#10 counter$count = 47999;
	#10 counter$count = 48000;
	#10 counter$count = 48001;
	#10 counter$count = 48002;
	#10 counter$count = 48003;
	#10 counter$count = 48004;
	#10 counter$count = 48005;
	#10 counter$count = 48006;
	#10 counter$count = 48007;
	#10 counter$count = 48008;
	#10 counter$count = 48009;
	#10 counter$count = 48010;
	#10 counter$count = 48011;
	#10 counter$count = 48012;
	#10 counter$count = 48013;
	#10 counter$count = 48014;
	#10 counter$count = 48015;
	#10 counter$count = 48016;
	#10 counter$count = 48017;
	#10 counter$count = 48018;
	#10 counter$count = 48019;
	#10 counter$count = 48020;
	#10 counter$count = 48021;
	#10 counter$count = 48022;
	#10 counter$count = 48023;
	#10 counter$count = 48024;
	#10 counter$count = 48025;
	#10 counter$count = 48026;
	#10 counter$count = 48027;
	#10 counter$count = 48028;
	#10 counter$count = 48029;
	#10 counter$count = 48030;
	#10 counter$count = 48031;
	#10 counter$count = 48032;
	#10 counter$count = 48033;
	#10 counter$count = 48034;
	#10 counter$count = 48035;
	#10 counter$count = 48036;
	#10 counter$count = 48037;
	#10 counter$count = 48038;
	#10 counter$count = 48039;
	#10 counter$count = 48040;
	#10 counter$count = 48041;
	#10 counter$count = 48042;
	#10 counter$count = 48043;
	#10 counter$count = 48044;
	#10 counter$count = 48045;
	#10 counter$count = 48046;
	#10 counter$count = 48047;
	#10 counter$count = 48048;
	#10 counter$count = 48049;
	#10 counter$count = 48050;
	#10 counter$count = 48051;
	#10 counter$count = 48052;
	#10 counter$count = 48053;
	#10 counter$count = 48054;
	#10 counter$count = 48055;
	#10 counter$count = 48056;
	#10 counter$count = 48057;
	#10 counter$count = 48058;
	#10 counter$count = 48059;
	#10 counter$count = 48060;
	#10 counter$count = 48061;
	#10 counter$count = 48062;
	#10 counter$count = 48063;
	#10 counter$count = 48064;
	#10 counter$count = 48065;
	#10 counter$count = 48066;
	#10 counter$count = 48067;
	#10 counter$count = 48068;
	#10 counter$count = 48069;
	#10 counter$count = 48070;
	#10 counter$count = 48071;
	#10 counter$count = 48072;
	#10 counter$count = 48073;
	#10 counter$count = 48074;
	#10 counter$count = 48075;
	#10 counter$count = 48076;
	#10 counter$count = 48077;
	#10 counter$count = 48078;
	#10 counter$count = 48079;
	#10 counter$count = 48080;
	#10 counter$count = 48081;
	#10 counter$count = 48082;
	#10 counter$count = 48083;
	#10 counter$count = 48084;
	#10 counter$count = 48085;
	#10 counter$count = 48086;
	#10 counter$count = 48087;
	#10 counter$count = 48088;
	#10 counter$count = 48089;
	#10 counter$count = 48090;
	#10 counter$count = 48091;
	#10 counter$count = 48092;
	#10 counter$count = 48093;
	#10 counter$count = 48094;
	#10 counter$count = 48095;
	#10 counter$count = 48096;
	#10 counter$count = 48097;
	#10 counter$count = 48098;
	#10 counter$count = 48099;
	#10 counter$count = 48100;
	#10 counter$count = 48101;
	#10 counter$count = 48102;
	#10 counter$count = 48103;
	#10 counter$count = 48104;
	#10 counter$count = 48105;
	#10 counter$count = 48106;
	#10 counter$count = 48107;
	#10 counter$count = 48108;
	#10 counter$count = 48109;
	#10 counter$count = 48110;
	#10 counter$count = 48111;
	#10 counter$count = 48112;
	#10 counter$count = 48113;
	#10 counter$count = 48114;
	#10 counter$count = 48115;
	#10 counter$count = 48116;
	#10 counter$count = 48117;
	#10 counter$count = 48118;
	#10 counter$count = 48119;
	#10 counter$count = 48120;
	#10 counter$count = 48121;
	#10 counter$count = 48122;
	#10 counter$count = 48123;
	#10 counter$count = 48124;
	#10 counter$count = 48125;
	#10 counter$count = 48126;
	#10 counter$count = 48127;
	#10 counter$count = 48128;
	#10 counter$count = 48129;
	#10 counter$count = 48130;
	#10 counter$count = 48131;
	#10 counter$count = 48132;
	#10 counter$count = 48133;
	#10 counter$count = 48134;
	#10 counter$count = 48135;
	#10 counter$count = 48136;
	#10 counter$count = 48137;
	#10 counter$count = 48138;
	#10 counter$count = 48139;
	#10 counter$count = 48140;
	#10 counter$count = 48141;
	#10 counter$count = 48142;
	#10 counter$count = 48143;
	#10 counter$count = 48144;
	#10 counter$count = 48145;
	#10 counter$count = 48146;
	#10 counter$count = 48147;
	#10 counter$count = 48148;
	#10 counter$count = 48149;
	#10 counter$count = 48150;
	#10 counter$count = 48151;
	#10 counter$count = 48152;
	#10 counter$count = 48153;
	#10 counter$count = 48154;
	#10 counter$count = 48155;
	#10 counter$count = 48156;
	#10 counter$count = 48157;
	#10 counter$count = 48158;
	#10 counter$count = 48159;
	#10 counter$count = 48160;
	#10 counter$count = 48161;
	#10 counter$count = 48162;
	#10 counter$count = 48163;
	#10 counter$count = 48164;
	#10 counter$count = 48165;
	#10 counter$count = 48166;
	#10 counter$count = 48167;
	#10 counter$count = 48168;
	#10 counter$count = 48169;
	#10 counter$count = 48170;
	#10 counter$count = 48171;
	#10 counter$count = 48172;
	#10 counter$count = 48173;
	#10 counter$count = 48174;
	#10 counter$count = 48175;
	#10 counter$count = 48176;
	#10 counter$count = 48177;
	#10 counter$count = 48178;
	#10 counter$count = 48179;
	#10 counter$count = 48180;
	#10 counter$count = 48181;
	#10 counter$count = 48182;
	#10 counter$count = 48183;
	#10 counter$count = 48184;
	#10 counter$count = 48185;
	#10 counter$count = 48186;
	#10 counter$count = 48187;
	#10 counter$count = 48188;
	#10 counter$count = 48189;
	#10 counter$count = 48190;
	#10 counter$count = 48191;
	#10 counter$count = 48192;
	#10 counter$count = 48193;
	#10 counter$count = 48194;
	#10 counter$count = 48195;
	#10 counter$count = 48196;
	#10 counter$count = 48197;
	#10 counter$count = 48198;
	#10 counter$count = 48199;
	#10 counter$count = 48200;
	#10 counter$count = 48201;
	#10 counter$count = 48202;
	#10 counter$count = 48203;
	#10 counter$count = 48204;
	#10 counter$count = 48205;
	#10 counter$count = 48206;
	#10 counter$count = 48207;
	#10 counter$count = 48208;
	#10 counter$count = 48209;
	#10 counter$count = 48210;
	#10 counter$count = 48211;
	#10 counter$count = 48212;
	#10 counter$count = 48213;
	#10 counter$count = 48214;
	#10 counter$count = 48215;
	#10 counter$count = 48216;
	#10 counter$count = 48217;
	#10 counter$count = 48218;
	#10 counter$count = 48219;
	#10 counter$count = 48220;
	#10 counter$count = 48221;
	#10 counter$count = 48222;
	#10 counter$count = 48223;
	#10 counter$count = 48224;
	#10 counter$count = 48225;
	#10 counter$count = 48226;
	#10 counter$count = 48227;
	#10 counter$count = 48228;
	#10 counter$count = 48229;
	#10 counter$count = 48230;
	#10 counter$count = 48231;
	#10 counter$count = 48232;
	#10 counter$count = 48233;
	#10 counter$count = 48234;
	#10 counter$count = 48235;
	#10 counter$count = 48236;
	#10 counter$count = 48237;
	#10 counter$count = 48238;
	#10 counter$count = 48239;
	#10 counter$count = 48240;
	#10 counter$count = 48241;
	#10 counter$count = 48242;
	#10 counter$count = 48243;
	#10 counter$count = 48244;
	#10 counter$count = 48245;
	#10 counter$count = 48246;
	#10 counter$count = 48247;
	#10 counter$count = 48248;
	#10 counter$count = 48249;
	#10 counter$count = 48250;
	#10 counter$count = 48251;
	#10 counter$count = 48252;
	#10 counter$count = 48253;
	#10 counter$count = 48254;
	#10 counter$count = 48255;
	#10 counter$count = 48256;
	#10 counter$count = 48257;
	#10 counter$count = 48258;
	#10 counter$count = 48259;
	#10 counter$count = 48260;
	#10 counter$count = 48261;
	#10 counter$count = 48262;
	#10 counter$count = 48263;
	#10 counter$count = 48264;
	#10 counter$count = 48265;
	#10 counter$count = 48266;
	#10 counter$count = 48267;
	#10 counter$count = 48268;
	#10 counter$count = 48269;
	#10 counter$count = 48270;
	#10 counter$count = 48271;
	#10 counter$count = 48272;
	#10 counter$count = 48273;
	#10 counter$count = 48274;
	#10 counter$count = 48275;
	#10 counter$count = 48276;
	#10 counter$count = 48277;
	#10 counter$count = 48278;
	#10 counter$count = 48279;
	#10 counter$count = 48280;
	#10 counter$count = 48281;
	#10 counter$count = 48282;
	#10 counter$count = 48283;
	#10 counter$count = 48284;
	#10 counter$count = 48285;
	#10 counter$count = 48286;
	#10 counter$count = 48287;
	#10 counter$count = 48288;
	#10 counter$count = 48289;
	#10 counter$count = 48290;
	#10 counter$count = 48291;
	#10 counter$count = 48292;
	#10 counter$count = 48293;
	#10 counter$count = 48294;
	#10 counter$count = 48295;
	#10 counter$count = 48296;
	#10 counter$count = 48297;
	#10 counter$count = 48298;
	#10 counter$count = 48299;
	#10 counter$count = 48300;
	#10 counter$count = 48301;
	#10 counter$count = 48302;
	#10 counter$count = 48303;
	#10 counter$count = 48304;
	#10 counter$count = 48305;
	#10 counter$count = 48306;
	#10 counter$count = 48307;
	#10 counter$count = 48308;
	#10 counter$count = 48309;
	#10 counter$count = 48310;
	#10 counter$count = 48311;
	#10 counter$count = 48312;
	#10 counter$count = 48313;
	#10 counter$count = 48314;
	#10 counter$count = 48315;
	#10 counter$count = 48316;
	#10 counter$count = 48317;
	#10 counter$count = 48318;
	#10 counter$count = 48319;
	#10 counter$count = 48320;
	#10 counter$count = 48321;
	#10 counter$count = 48322;
	#10 counter$count = 48323;
	#10 counter$count = 48324;
	#10 counter$count = 48325;
	#10 counter$count = 48326;
	#10 counter$count = 48327;
	#10 counter$count = 48328;
	#10 counter$count = 48329;
	#10 counter$count = 48330;
	#10 counter$count = 48331;
	#10 counter$count = 48332;
	#10 counter$count = 48333;
	#10 counter$count = 48334;
	#10 counter$count = 48335;
	#10 counter$count = 48336;
	#10 counter$count = 48337;
	#10 counter$count = 48338;
	#10 counter$count = 48339;
	#10 counter$count = 48340;
	#10 counter$count = 48341;
	#10 counter$count = 48342;
	#10 counter$count = 48343;
	#10 counter$count = 48344;
	#10 counter$count = 48345;
	#10 counter$count = 48346;
	#10 counter$count = 48347;
	#10 counter$count = 48348;
	#10 counter$count = 48349;
	#10 counter$count = 48350;
	#10 counter$count = 48351;
	#10 counter$count = 48352;
	#10 counter$count = 48353;
	#10 counter$count = 48354;
	#10 counter$count = 48355;
	#10 counter$count = 48356;
	#10 counter$count = 48357;
	#10 counter$count = 48358;
	#10 counter$count = 48359;
	#10 counter$count = 48360;
	#10 counter$count = 48361;
	#10 counter$count = 48362;
	#10 counter$count = 48363;
	#10 counter$count = 48364;
	#10 counter$count = 48365;
	#10 counter$count = 48366;
	#10 counter$count = 48367;
	#10 counter$count = 48368;
	#10 counter$count = 48369;
	#10 counter$count = 48370;
	#10 counter$count = 48371;
	#10 counter$count = 48372;
	#10 counter$count = 48373;
	#10 counter$count = 48374;
	#10 counter$count = 48375;
	#10 counter$count = 48376;
	#10 counter$count = 48377;
	#10 counter$count = 48378;
	#10 counter$count = 48379;
	#10 counter$count = 48380;
	#10 counter$count = 48381;
	#10 counter$count = 48382;
	#10 counter$count = 48383;
	#10 counter$count = 48384;
	#10 counter$count = 48385;
	#10 counter$count = 48386;
	#10 counter$count = 48387;
	#10 counter$count = 48388;
	#10 counter$count = 48389;
	#10 counter$count = 48390;
	#10 counter$count = 48391;
	#10 counter$count = 48392;
	#10 counter$count = 48393;
	#10 counter$count = 48394;
	#10 counter$count = 48395;
	#10 counter$count = 48396;
	#10 counter$count = 48397;
	#10 counter$count = 48398;
	#10 counter$count = 48399;
	#10 counter$count = 48400;
	#10 counter$count = 48401;
	#10 counter$count = 48402;
	#10 counter$count = 48403;
	#10 counter$count = 48404;
	#10 counter$count = 48405;
	#10 counter$count = 48406;
	#10 counter$count = 48407;
	#10 counter$count = 48408;
	#10 counter$count = 48409;
	#10 counter$count = 48410;
	#10 counter$count = 48411;
	#10 counter$count = 48412;
	#10 counter$count = 48413;
	#10 counter$count = 48414;
	#10 counter$count = 48415;
	#10 counter$count = 48416;
	#10 counter$count = 48417;
	#10 counter$count = 48418;
	#10 counter$count = 48419;
	#10 counter$count = 48420;
	#10 counter$count = 48421;
	#10 counter$count = 48422;
	#10 counter$count = 48423;
	#10 counter$count = 48424;
	#10 counter$count = 48425;
	#10 counter$count = 48426;
	#10 counter$count = 48427;
	#10 counter$count = 48428;
	#10 counter$count = 48429;
	#10 counter$count = 48430;
	#10 counter$count = 48431;
	#10 counter$count = 48432;
	#10 counter$count = 48433;
	#10 counter$count = 48434;
	#10 counter$count = 48435;
	#10 counter$count = 48436;
	#10 counter$count = 48437;
	#10 counter$count = 48438;
	#10 counter$count = 48439;
	#10 counter$count = 48440;
	#10 counter$count = 48441;
	#10 counter$count = 48442;
	#10 counter$count = 48443;
	#10 counter$count = 48444;
	#10 counter$count = 48445;
	#10 counter$count = 48446;
	#10 counter$count = 48447;
	#10 counter$count = 48448;
	#10 counter$count = 48449;
	#10 counter$count = 48450;
	#10 counter$count = 48451;
	#10 counter$count = 48452;
	#10 counter$count = 48453;
	#10 counter$count = 48454;
	#10 counter$count = 48455;
	#10 counter$count = 48456;
	#10 counter$count = 48457;
	#10 counter$count = 48458;
	#10 counter$count = 48459;
	#10 counter$count = 48460;
	#10 counter$count = 48461;
	#10 counter$count = 48462;
	#10 counter$count = 48463;
	#10 counter$count = 48464;
	#10 counter$count = 48465;
	#10 counter$count = 48466;
	#10 counter$count = 48467;
	#10 counter$count = 48468;
	#10 counter$count = 48469;
	#10 counter$count = 48470;
	#10 counter$count = 48471;
	#10 counter$count = 48472;
	#10 counter$count = 48473;
	#10 counter$count = 48474;
	#10 counter$count = 48475;
	#10 counter$count = 48476;
	#10 counter$count = 48477;
	#10 counter$count = 48478;
	#10 counter$count = 48479;
	#10 counter$count = 48480;
	#10 counter$count = 48481;
	#10 counter$count = 48482;
	#10 counter$count = 48483;
	#10 counter$count = 48484;
	#10 counter$count = 48485;
	#10 counter$count = 48486;
	#10 counter$count = 48487;
	#10 counter$count = 48488;
	#10 counter$count = 48489;
	#10 counter$count = 48490;
	#10 counter$count = 48491;
	#10 counter$count = 48492;
	#10 counter$count = 48493;
	#10 counter$count = 48494;
	#10 counter$count = 48495;
	#10 counter$count = 48496;
	#10 counter$count = 48497;
	#10 counter$count = 48498;
	#10 counter$count = 48499;
	#10 counter$count = 48500;
	#10 counter$count = 48501;
	#10 counter$count = 48502;
	#10 counter$count = 48503;
	#10 counter$count = 48504;
	#10 counter$count = 48505;
	#10 counter$count = 48506;
	#10 counter$count = 48507;
	#10 counter$count = 48508;
	#10 counter$count = 48509;
	#10 counter$count = 48510;
	#10 counter$count = 48511;
	#10 counter$count = 48512;
	#10 counter$count = 48513;
	#10 counter$count = 48514;
	#10 counter$count = 48515;
	#10 counter$count = 48516;
	#10 counter$count = 48517;
	#10 counter$count = 48518;
	#10 counter$count = 48519;
	#10 counter$count = 48520;
	#10 counter$count = 48521;
	#10 counter$count = 48522;
	#10 counter$count = 48523;
	#10 counter$count = 48524;
	#10 counter$count = 48525;
	#10 counter$count = 48526;
	#10 counter$count = 48527;
	#10 counter$count = 48528;
	#10 counter$count = 48529;
	#10 counter$count = 48530;
	#10 counter$count = 48531;
	#10 counter$count = 48532;
	#10 counter$count = 48533;
	#10 counter$count = 48534;
	#10 counter$count = 48535;
	#10 counter$count = 48536;
	#10 counter$count = 48537;
	#10 counter$count = 48538;
	#10 counter$count = 48539;
	#10 counter$count = 48540;
	#10 counter$count = 48541;
	#10 counter$count = 48542;
	#10 counter$count = 48543;
	#10 counter$count = 48544;
	#10 counter$count = 48545;
	#10 counter$count = 48546;
	#10 counter$count = 48547;
	#10 counter$count = 48548;
	#10 counter$count = 48549;
	#10 counter$count = 48550;
	#10 counter$count = 48551;
	#10 counter$count = 48552;
	#10 counter$count = 48553;
	#10 counter$count = 48554;
	#10 counter$count = 48555;
	#10 counter$count = 48556;
	#10 counter$count = 48557;
	#10 counter$count = 48558;
	#10 counter$count = 48559;
	#10 counter$count = 48560;
	#10 counter$count = 48561;
	#10 counter$count = 48562;
	#10 counter$count = 48563;
	#10 counter$count = 48564;
	#10 counter$count = 48565;
	#10 counter$count = 48566;
	#10 counter$count = 48567;
	#10 counter$count = 48568;
	#10 counter$count = 48569;
	#10 counter$count = 48570;
	#10 counter$count = 48571;
	#10 counter$count = 48572;
	#10 counter$count = 48573;
	#10 counter$count = 48574;
	#10 counter$count = 48575;
	#10 counter$count = 48576;
	#10 counter$count = 48577;
	#10 counter$count = 48578;
	#10 counter$count = 48579;
	#10 counter$count = 48580;
	#10 counter$count = 48581;
	#10 counter$count = 48582;
	#10 counter$count = 48583;
	#10 counter$count = 48584;
	#10 counter$count = 48585;
	#10 counter$count = 48586;
	#10 counter$count = 48587;
	#10 counter$count = 48588;
	#10 counter$count = 48589;
	#10 counter$count = 48590;
	#10 counter$count = 48591;
	#10 counter$count = 48592;
	#10 counter$count = 48593;
	#10 counter$count = 48594;
	#10 counter$count = 48595;
	#10 counter$count = 48596;
	#10 counter$count = 48597;
	#10 counter$count = 48598;
	#10 counter$count = 48599;
	#10 counter$count = 48600;
	#10 counter$count = 48601;
	#10 counter$count = 48602;
	#10 counter$count = 48603;
	#10 counter$count = 48604;
	#10 counter$count = 48605;
	#10 counter$count = 48606;
	#10 counter$count = 48607;
	#10 counter$count = 48608;
	#10 counter$count = 48609;
	#10 counter$count = 48610;
	#10 counter$count = 48611;
	#10 counter$count = 48612;
	#10 counter$count = 48613;
	#10 counter$count = 48614;
	#10 counter$count = 48615;
	#10 counter$count = 48616;
	#10 counter$count = 48617;
	#10 counter$count = 48618;
	#10 counter$count = 48619;
	#10 counter$count = 48620;
	#10 counter$count = 48621;
	#10 counter$count = 48622;
	#10 counter$count = 48623;
	#10 counter$count = 48624;
	#10 counter$count = 48625;
	#10 counter$count = 48626;
	#10 counter$count = 48627;
	#10 counter$count = 48628;
	#10 counter$count = 48629;
	#10 counter$count = 48630;
	#10 counter$count = 48631;
	#10 counter$count = 48632;
	#10 counter$count = 48633;
	#10 counter$count = 48634;
	#10 counter$count = 48635;
	#10 counter$count = 48636;
	#10 counter$count = 48637;
	#10 counter$count = 48638;
	#10 counter$count = 48639;
	#10 counter$count = 48640;
	#10 counter$count = 48641;
	#10 counter$count = 48642;
	#10 counter$count = 48643;
	#10 counter$count = 48644;
	#10 counter$count = 48645;
	#10 counter$count = 48646;
	#10 counter$count = 48647;
	#10 counter$count = 48648;
	#10 counter$count = 48649;
	#10 counter$count = 48650;
	#10 counter$count = 48651;
	#10 counter$count = 48652;
	#10 counter$count = 48653;
	#10 counter$count = 48654;
	#10 counter$count = 48655;
	#10 counter$count = 48656;
	#10 counter$count = 48657;
	#10 counter$count = 48658;
	#10 counter$count = 48659;
	#10 counter$count = 48660;
	#10 counter$count = 48661;
	#10 counter$count = 48662;
	#10 counter$count = 48663;
	#10 counter$count = 48664;
	#10 counter$count = 48665;
	#10 counter$count = 48666;
	#10 counter$count = 48667;
	#10 counter$count = 48668;
	#10 counter$count = 48669;
	#10 counter$count = 48670;
	#10 counter$count = 48671;
	#10 counter$count = 48672;
	#10 counter$count = 48673;
	#10 counter$count = 48674;
	#10 counter$count = 48675;
	#10 counter$count = 48676;
	#10 counter$count = 48677;
	#10 counter$count = 48678;
	#10 counter$count = 48679;
	#10 counter$count = 48680;
	#10 counter$count = 48681;
	#10 counter$count = 48682;
	#10 counter$count = 48683;
	#10 counter$count = 48684;
	#10 counter$count = 48685;
	#10 counter$count = 48686;
	#10 counter$count = 48687;
	#10 counter$count = 48688;
	#10 counter$count = 48689;
	#10 counter$count = 48690;
	#10 counter$count = 48691;
	#10 counter$count = 48692;
	#10 counter$count = 48693;
	#10 counter$count = 48694;
	#10 counter$count = 48695;
	#10 counter$count = 48696;
	#10 counter$count = 48697;
	#10 counter$count = 48698;
	#10 counter$count = 48699;
	#10 counter$count = 48700;
	#10 counter$count = 48701;
	#10 counter$count = 48702;
	#10 counter$count = 48703;
	#10 counter$count = 48704;
	#10 counter$count = 48705;
	#10 counter$count = 48706;
	#10 counter$count = 48707;
	#10 counter$count = 48708;
	#10 counter$count = 48709;
	#10 counter$count = 48710;
	#10 counter$count = 48711;
	#10 counter$count = 48712;
	#10 counter$count = 48713;
	#10 counter$count = 48714;
	#10 counter$count = 48715;
	#10 counter$count = 48716;
	#10 counter$count = 48717;
	#10 counter$count = 48718;
	#10 counter$count = 48719;
	#10 counter$count = 48720;
	#10 counter$count = 48721;
	#10 counter$count = 48722;
	#10 counter$count = 48723;
	#10 counter$count = 48724;
	#10 counter$count = 48725;
	#10 counter$count = 48726;
	#10 counter$count = 48727;
	#10 counter$count = 48728;
	#10 counter$count = 48729;
	#10 counter$count = 48730;
	#10 counter$count = 48731;
	#10 counter$count = 48732;
	#10 counter$count = 48733;
	#10 counter$count = 48734;
	#10 counter$count = 48735;
	#10 counter$count = 48736;
	#10 counter$count = 48737;
	#10 counter$count = 48738;
	#10 counter$count = 48739;
	#10 counter$count = 48740;
	#10 counter$count = 48741;
	#10 counter$count = 48742;
	#10 counter$count = 48743;
	#10 counter$count = 48744;
	#10 counter$count = 48745;
	#10 counter$count = 48746;
	#10 counter$count = 48747;
	#10 counter$count = 48748;
	#10 counter$count = 48749;
	#10 counter$count = 48750;
	#10 counter$count = 48751;
	#10 counter$count = 48752;
	#10 counter$count = 48753;
	#10 counter$count = 48754;
	#10 counter$count = 48755;
	#10 counter$count = 48756;
	#10 counter$count = 48757;
	#10 counter$count = 48758;
	#10 counter$count = 48759;
	#10 counter$count = 48760;
	#10 counter$count = 48761;
	#10 counter$count = 48762;
	#10 counter$count = 48763;
	#10 counter$count = 48764;
	#10 counter$count = 48765;
	#10 counter$count = 48766;
	#10 counter$count = 48767;
	#10 counter$count = 48768;
	#10 counter$count = 48769;
	#10 counter$count = 48770;
	#10 counter$count = 48771;
	#10 counter$count = 48772;
	#10 counter$count = 48773;
	#10 counter$count = 48774;
	#10 counter$count = 48775;
	#10 counter$count = 48776;
	#10 counter$count = 48777;
	#10 counter$count = 48778;
	#10 counter$count = 48779;
	#10 counter$count = 48780;
	#10 counter$count = 48781;
	#10 counter$count = 48782;
	#10 counter$count = 48783;
	#10 counter$count = 48784;
	#10 counter$count = 48785;
	#10 counter$count = 48786;
	#10 counter$count = 48787;
	#10 counter$count = 48788;
	#10 counter$count = 48789;
	#10 counter$count = 48790;
	#10 counter$count = 48791;
	#10 counter$count = 48792;
	#10 counter$count = 48793;
	#10 counter$count = 48794;
	#10 counter$count = 48795;
	#10 counter$count = 48796;
	#10 counter$count = 48797;
	#10 counter$count = 48798;
	#10 counter$count = 48799;
	#10 counter$count = 48800;
	#10 counter$count = 48801;
	#10 counter$count = 48802;
	#10 counter$count = 48803;
	#10 counter$count = 48804;
	#10 counter$count = 48805;
	#10 counter$count = 48806;
	#10 counter$count = 48807;
	#10 counter$count = 48808;
	#10 counter$count = 48809;
	#10 counter$count = 48810;
	#10 counter$count = 48811;
	#10 counter$count = 48812;
	#10 counter$count = 48813;
	#10 counter$count = 48814;
	#10 counter$count = 48815;
	#10 counter$count = 48816;
	#10 counter$count = 48817;
	#10 counter$count = 48818;
	#10 counter$count = 48819;
	#10 counter$count = 48820;
	#10 counter$count = 48821;
	#10 counter$count = 48822;
	#10 counter$count = 48823;
	#10 counter$count = 48824;
	#10 counter$count = 48825;
	#10 counter$count = 48826;
	#10 counter$count = 48827;
	#10 counter$count = 48828;
	#10 counter$count = 48829;
	#10 counter$count = 48830;
	#10 counter$count = 48831;
	#10 counter$count = 48832;
	#10 counter$count = 48833;
	#10 counter$count = 48834;
	#10 counter$count = 48835;
	#10 counter$count = 48836;
	#10 counter$count = 48837;
	#10 counter$count = 48838;
	#10 counter$count = 48839;
	#10 counter$count = 48840;
	#10 counter$count = 48841;
	#10 counter$count = 48842;
	#10 counter$count = 48843;
	#10 counter$count = 48844;
	#10 counter$count = 48845;
	#10 counter$count = 48846;
	#10 counter$count = 48847;
	#10 counter$count = 48848;
	#10 counter$count = 48849;
	#10 counter$count = 48850;
	#10 counter$count = 48851;
	#10 counter$count = 48852;
	#10 counter$count = 48853;
	#10 counter$count = 48854;
	#10 counter$count = 48855;
	#10 counter$count = 48856;
	#10 counter$count = 48857;
	#10 counter$count = 48858;
	#10 counter$count = 48859;
	#10 counter$count = 48860;
	#10 counter$count = 48861;
	#10 counter$count = 48862;
	#10 counter$count = 48863;
	#10 counter$count = 48864;
	#10 counter$count = 48865;
	#10 counter$count = 48866;
	#10 counter$count = 48867;
	#10 counter$count = 48868;
	#10 counter$count = 48869;
	#10 counter$count = 48870;
	#10 counter$count = 48871;
	#10 counter$count = 48872;
	#10 counter$count = 48873;
	#10 counter$count = 48874;
	#10 counter$count = 48875;
	#10 counter$count = 48876;
	#10 counter$count = 48877;
	#10 counter$count = 48878;
	#10 counter$count = 48879;
	#10 counter$count = 48880;
	#10 counter$count = 48881;
	#10 counter$count = 48882;
	#10 counter$count = 48883;
	#10 counter$count = 48884;
	#10 counter$count = 48885;
	#10 counter$count = 48886;
	#10 counter$count = 48887;
	#10 counter$count = 48888;
	#10 counter$count = 48889;
	#10 counter$count = 48890;
	#10 counter$count = 48891;
	#10 counter$count = 48892;
	#10 counter$count = 48893;
	#10 counter$count = 48894;
	#10 counter$count = 48895;
	#10 counter$count = 48896;
	#10 counter$count = 48897;
	#10 counter$count = 48898;
	#10 counter$count = 48899;
	#10 counter$count = 48900;
	#10 counter$count = 48901;
	#10 counter$count = 48902;
	#10 counter$count = 48903;
	#10 counter$count = 48904;
	#10 counter$count = 48905;
	#10 counter$count = 48906;
	#10 counter$count = 48907;
	#10 counter$count = 48908;
	#10 counter$count = 48909;
	#10 counter$count = 48910;
	#10 counter$count = 48911;
	#10 counter$count = 48912;
	#10 counter$count = 48913;
	#10 counter$count = 48914;
	#10 counter$count = 48915;
	#10 counter$count = 48916;
	#10 counter$count = 48917;
	#10 counter$count = 48918;
	#10 counter$count = 48919;
	#10 counter$count = 48920;
	#10 counter$count = 48921;
	#10 counter$count = 48922;
	#10 counter$count = 48923;
	#10 counter$count = 48924;
	#10 counter$count = 48925;
	#10 counter$count = 48926;
	#10 counter$count = 48927;
	#10 counter$count = 48928;
	#10 counter$count = 48929;
	#10 counter$count = 48930;
	#10 counter$count = 48931;
	#10 counter$count = 48932;
	#10 counter$count = 48933;
	#10 counter$count = 48934;
	#10 counter$count = 48935;
	#10 counter$count = 48936;
	#10 counter$count = 48937;
	#10 counter$count = 48938;
	#10 counter$count = 48939;
	#10 counter$count = 48940;
	#10 counter$count = 48941;
	#10 counter$count = 48942;
	#10 counter$count = 48943;
	#10 counter$count = 48944;
	#10 counter$count = 48945;
	#10 counter$count = 48946;
	#10 counter$count = 48947;
	#10 counter$count = 48948;
	#10 counter$count = 48949;
	#10 counter$count = 48950;
	#10 counter$count = 48951;
	#10 counter$count = 48952;
	#10 counter$count = 48953;
	#10 counter$count = 48954;
	#10 counter$count = 48955;
	#10 counter$count = 48956;
	#10 counter$count = 48957;
	#10 counter$count = 48958;
	#10 counter$count = 48959;
	#10 counter$count = 48960;
	#10 counter$count = 48961;
	#10 counter$count = 48962;
	#10 counter$count = 48963;
	#10 counter$count = 48964;
	#10 counter$count = 48965;
	#10 counter$count = 48966;
	#10 counter$count = 48967;
	#10 counter$count = 48968;
	#10 counter$count = 48969;
	#10 counter$count = 48970;
	#10 counter$count = 48971;
	#10 counter$count = 48972;
	#10 counter$count = 48973;
	#10 counter$count = 48974;
	#10 counter$count = 48975;
	#10 counter$count = 48976;
	#10 counter$count = 48977;
	#10 counter$count = 48978;
	#10 counter$count = 48979;
	#10 counter$count = 48980;
	#10 counter$count = 48981;
	#10 counter$count = 48982;
	#10 counter$count = 48983;
	#10 counter$count = 48984;
	#10 counter$count = 48985;
	#10 counter$count = 48986;
	#10 counter$count = 48987;
	#10 counter$count = 48988;
	#10 counter$count = 48989;
	#10 counter$count = 48990;
	#10 counter$count = 48991;
	#10 counter$count = 48992;
	#10 counter$count = 48993;
	#10 counter$count = 48994;
	#10 counter$count = 48995;
	#10 counter$count = 48996;
	#10 counter$count = 48997;
	#10 counter$count = 48998;
	#10 counter$count = 48999;
	#10 counter$count = 49000;
	#10 counter$count = 49001;
	#10 counter$count = 49002;
	#10 counter$count = 49003;
	#10 counter$count = 49004;
	#10 counter$count = 49005;
	#10 counter$count = 49006;
	#10 counter$count = 49007;
	#10 counter$count = 49008;
	#10 counter$count = 49009;
	#10 counter$count = 49010;
	#10 counter$count = 49011;
	#10 counter$count = 49012;
	#10 counter$count = 49013;
	#10 counter$count = 49014;
	#10 counter$count = 49015;
	#10 counter$count = 49016;
	#10 counter$count = 49017;
	#10 counter$count = 49018;
	#10 counter$count = 49019;
	#10 counter$count = 49020;
	#10 counter$count = 49021;
	#10 counter$count = 49022;
	#10 counter$count = 49023;
	#10 counter$count = 49024;
	#10 counter$count = 49025;
	#10 counter$count = 49026;
	#10 counter$count = 49027;
	#10 counter$count = 49028;
	#10 counter$count = 49029;
	#10 counter$count = 49030;
	#10 counter$count = 49031;
	#10 counter$count = 49032;
	#10 counter$count = 49033;
	#10 counter$count = 49034;
	#10 counter$count = 49035;
	#10 counter$count = 49036;
	#10 counter$count = 49037;
	#10 counter$count = 49038;
	#10 counter$count = 49039;
	#10 counter$count = 49040;
	#10 counter$count = 49041;
	#10 counter$count = 49042;
	#10 counter$count = 49043;
	#10 counter$count = 49044;
	#10 counter$count = 49045;
	#10 counter$count = 49046;
	#10 counter$count = 49047;
	#10 counter$count = 49048;
	#10 counter$count = 49049;
	#10 counter$count = 49050;
	#10 counter$count = 49051;
	#10 counter$count = 49052;
	#10 counter$count = 49053;
	#10 counter$count = 49054;
	#10 counter$count = 49055;
	#10 counter$count = 49056;
	#10 counter$count = 49057;
	#10 counter$count = 49058;
	#10 counter$count = 49059;
	#10 counter$count = 49060;
	#10 counter$count = 49061;
	#10 counter$count = 49062;
	#10 counter$count = 49063;
	#10 counter$count = 49064;
	#10 counter$count = 49065;
	#10 counter$count = 49066;
	#10 counter$count = 49067;
	#10 counter$count = 49068;
	#10 counter$count = 49069;
	#10 counter$count = 49070;
	#10 counter$count = 49071;
	#10 counter$count = 49072;
	#10 counter$count = 49073;
	#10 counter$count = 49074;
	#10 counter$count = 49075;
	#10 counter$count = 49076;
	#10 counter$count = 49077;
	#10 counter$count = 49078;
	#10 counter$count = 49079;
	#10 counter$count = 49080;
	#10 counter$count = 49081;
	#10 counter$count = 49082;
	#10 counter$count = 49083;
	#10 counter$count = 49084;
	#10 counter$count = 49085;
	#10 counter$count = 49086;
	#10 counter$count = 49087;
	#10 counter$count = 49088;
	#10 counter$count = 49089;
	#10 counter$count = 49090;
	#10 counter$count = 49091;
	#10 counter$count = 49092;
	#10 counter$count = 49093;
	#10 counter$count = 49094;
	#10 counter$count = 49095;
	#10 counter$count = 49096;
	#10 counter$count = 49097;
	#10 counter$count = 49098;
	#10 counter$count = 49099;
	#10 counter$count = 49100;
	#10 counter$count = 49101;
	#10 counter$count = 49102;
	#10 counter$count = 49103;
	#10 counter$count = 49104;
	#10 counter$count = 49105;
	#10 counter$count = 49106;
	#10 counter$count = 49107;
	#10 counter$count = 49108;
	#10 counter$count = 49109;
	#10 counter$count = 49110;
	#10 counter$count = 49111;
	#10 counter$count = 49112;
	#10 counter$count = 49113;
	#10 counter$count = 49114;
	#10 counter$count = 49115;
	#10 counter$count = 49116;
	#10 counter$count = 49117;
	#10 counter$count = 49118;
	#10 counter$count = 49119;
	#10 counter$count = 49120;
	#10 counter$count = 49121;
	#10 counter$count = 49122;
	#10 counter$count = 49123;
	#10 counter$count = 49124;
	#10 counter$count = 49125;
	#10 counter$count = 49126;
	#10 counter$count = 49127;
	#10 counter$count = 49128;
	#10 counter$count = 49129;
	#10 counter$count = 49130;
	#10 counter$count = 49131;
	#10 counter$count = 49132;
	#10 counter$count = 49133;
	#10 counter$count = 49134;
	#10 counter$count = 49135;
	#10 counter$count = 49136;
	#10 counter$count = 49137;
	#10 counter$count = 49138;
	#10 counter$count = 49139;
	#10 counter$count = 49140;
	#10 counter$count = 49141;
	#10 counter$count = 49142;
	#10 counter$count = 49143;
	#10 counter$count = 49144;
	#10 counter$count = 49145;
	#10 counter$count = 49146;
	#10 counter$count = 49147;
	#10 counter$count = 49148;
	#10 counter$count = 49149;
	#10 counter$count = 49150;
	#10 counter$count = 49151;
	#10 counter$count = 49152;
	#10 counter$count = 49153;
	#10 counter$count = 49154;
	#10 counter$count = 49155;
	#10 counter$count = 49156;
	#10 counter$count = 49157;
	#10 counter$count = 49158;
	#10 counter$count = 49159;
	#10 counter$count = 49160;
	#10 counter$count = 49161;
	#10 counter$count = 49162;
	#10 counter$count = 49163;
	#10 counter$count = 49164;
	#10 counter$count = 49165;
	#10 counter$count = 49166;
	#10 counter$count = 49167;
	#10 counter$count = 49168;
	#10 counter$count = 49169;
	#10 counter$count = 49170;
	#10 counter$count = 49171;
	#10 counter$count = 49172;
	#10 counter$count = 49173;
	#10 counter$count = 49174;
	#10 counter$count = 49175;
	#10 counter$count = 49176;
	#10 counter$count = 49177;
	#10 counter$count = 49178;
	#10 counter$count = 49179;
	#10 counter$count = 49180;
	#10 counter$count = 49181;
	#10 counter$count = 49182;
	#10 counter$count = 49183;
	#10 counter$count = 49184;
	#10 counter$count = 49185;
	#10 counter$count = 49186;
	#10 counter$count = 49187;
	#10 counter$count = 49188;
	#10 counter$count = 49189;
	#10 counter$count = 49190;
	#10 counter$count = 49191;
	#10 counter$count = 49192;
	#10 counter$count = 49193;
	#10 counter$count = 49194;
	#10 counter$count = 49195;
	#10 counter$count = 49196;
	#10 counter$count = 49197;
	#10 counter$count = 49198;
	#10 counter$count = 49199;
	#10 counter$count = 49200;
	#10 counter$count = 49201;
	#10 counter$count = 49202;
	#10 counter$count = 49203;
	#10 counter$count = 49204;
	#10 counter$count = 49205;
	#10 counter$count = 49206;
	#10 counter$count = 49207;
	#10 counter$count = 49208;
	#10 counter$count = 49209;
	#10 counter$count = 49210;
	#10 counter$count = 49211;
	#10 counter$count = 49212;
	#10 counter$count = 49213;
	#10 counter$count = 49214;
	#10 counter$count = 49215;
	#10 counter$count = 49216;
	#10 counter$count = 49217;
	#10 counter$count = 49218;
	#10 counter$count = 49219;
	#10 counter$count = 49220;
	#10 counter$count = 49221;
	#10 counter$count = 49222;
	#10 counter$count = 49223;
	#10 counter$count = 49224;
	#10 counter$count = 49225;
	#10 counter$count = 49226;
	#10 counter$count = 49227;
	#10 counter$count = 49228;
	#10 counter$count = 49229;
	#10 counter$count = 49230;
	#10 counter$count = 49231;
	#10 counter$count = 49232;
	#10 counter$count = 49233;
	#10 counter$count = 49234;
	#10 counter$count = 49235;
	#10 counter$count = 49236;
	#10 counter$count = 49237;
	#10 counter$count = 49238;
	#10 counter$count = 49239;
	#10 counter$count = 49240;
	#10 counter$count = 49241;
	#10 counter$count = 49242;
	#10 counter$count = 49243;
	#10 counter$count = 49244;
	#10 counter$count = 49245;
	#10 counter$count = 49246;
	#10 counter$count = 49247;
	#10 counter$count = 49248;
	#10 counter$count = 49249;
	#10 counter$count = 49250;
	#10 counter$count = 49251;
	#10 counter$count = 49252;
	#10 counter$count = 49253;
	#10 counter$count = 49254;
	#10 counter$count = 49255;
	#10 counter$count = 49256;
	#10 counter$count = 49257;
	#10 counter$count = 49258;
	#10 counter$count = 49259;
	#10 counter$count = 49260;
	#10 counter$count = 49261;
	#10 counter$count = 49262;
	#10 counter$count = 49263;
	#10 counter$count = 49264;
	#10 counter$count = 49265;
	#10 counter$count = 49266;
	#10 counter$count = 49267;
	#10 counter$count = 49268;
	#10 counter$count = 49269;
	#10 counter$count = 49270;
	#10 counter$count = 49271;
	#10 counter$count = 49272;
	#10 counter$count = 49273;
	#10 counter$count = 49274;
	#10 counter$count = 49275;
	#10 counter$count = 49276;
	#10 counter$count = 49277;
	#10 counter$count = 49278;
	#10 counter$count = 49279;
	#10 counter$count = 49280;
	#10 counter$count = 49281;
	#10 counter$count = 49282;
	#10 counter$count = 49283;
	#10 counter$count = 49284;
	#10 counter$count = 49285;
	#10 counter$count = 49286;
	#10 counter$count = 49287;
	#10 counter$count = 49288;
	#10 counter$count = 49289;
	#10 counter$count = 49290;
	#10 counter$count = 49291;
	#10 counter$count = 49292;
	#10 counter$count = 49293;
	#10 counter$count = 49294;
	#10 counter$count = 49295;
	#10 counter$count = 49296;
	#10 counter$count = 49297;
	#10 counter$count = 49298;
	#10 counter$count = 49299;
	#10 counter$count = 49300;
	#10 counter$count = 49301;
	#10 counter$count = 49302;
	#10 counter$count = 49303;
	#10 counter$count = 49304;
	#10 counter$count = 49305;
	#10 counter$count = 49306;
	#10 counter$count = 49307;
	#10 counter$count = 49308;
	#10 counter$count = 49309;
	#10 counter$count = 49310;
	#10 counter$count = 49311;
	#10 counter$count = 49312;
	#10 counter$count = 49313;
	#10 counter$count = 49314;
	#10 counter$count = 49315;
	#10 counter$count = 49316;
	#10 counter$count = 49317;
	#10 counter$count = 49318;
	#10 counter$count = 49319;
	#10 counter$count = 49320;
	#10 counter$count = 49321;
	#10 counter$count = 49322;
	#10 counter$count = 49323;
	#10 counter$count = 49324;
	#10 counter$count = 49325;
	#10 counter$count = 49326;
	#10 counter$count = 49327;
	#10 counter$count = 49328;
	#10 counter$count = 49329;
	#10 counter$count = 49330;
	#10 counter$count = 49331;
	#10 counter$count = 49332;
	#10 counter$count = 49333;
	#10 counter$count = 49334;
	#10 counter$count = 49335;
	#10 counter$count = 49336;
	#10 counter$count = 49337;
	#10 counter$count = 49338;
	#10 counter$count = 49339;
	#10 counter$count = 49340;
	#10 counter$count = 49341;
	#10 counter$count = 49342;
	#10 counter$count = 49343;
	#10 counter$count = 49344;
	#10 counter$count = 49345;
	#10 counter$count = 49346;
	#10 counter$count = 49347;
	#10 counter$count = 49348;
	#10 counter$count = 49349;
	#10 counter$count = 49350;
	#10 counter$count = 49351;
	#10 counter$count = 49352;
	#10 counter$count = 49353;
	#10 counter$count = 49354;
	#10 counter$count = 49355;
	#10 counter$count = 49356;
	#10 counter$count = 49357;
	#10 counter$count = 49358;
	#10 counter$count = 49359;
	#10 counter$count = 49360;
	#10 counter$count = 49361;
	#10 counter$count = 49362;
	#10 counter$count = 49363;
	#10 counter$count = 49364;
	#10 counter$count = 49365;
	#10 counter$count = 49366;
	#10 counter$count = 49367;
	#10 counter$count = 49368;
	#10 counter$count = 49369;
	#10 counter$count = 49370;
	#10 counter$count = 49371;
	#10 counter$count = 49372;
	#10 counter$count = 49373;
	#10 counter$count = 49374;
	#10 counter$count = 49375;
	#10 counter$count = 49376;
	#10 counter$count = 49377;
	#10 counter$count = 49378;
	#10 counter$count = 49379;
	#10 counter$count = 49380;
	#10 counter$count = 49381;
	#10 counter$count = 49382;
	#10 counter$count = 49383;
	#10 counter$count = 49384;
	#10 counter$count = 49385;
	#10 counter$count = 49386;
	#10 counter$count = 49387;
	#10 counter$count = 49388;
	#10 counter$count = 49389;
	#10 counter$count = 49390;
	#10 counter$count = 49391;
	#10 counter$count = 49392;
	#10 counter$count = 49393;
	#10 counter$count = 49394;
	#10 counter$count = 49395;
	#10 counter$count = 49396;
	#10 counter$count = 49397;
	#10 counter$count = 49398;
	#10 counter$count = 49399;
	#10 counter$count = 49400;
	#10 counter$count = 49401;
	#10 counter$count = 49402;
	#10 counter$count = 49403;
	#10 counter$count = 49404;
	#10 counter$count = 49405;
	#10 counter$count = 49406;
	#10 counter$count = 49407;
	#10 counter$count = 49408;
	#10 counter$count = 49409;
	#10 counter$count = 49410;
	#10 counter$count = 49411;
	#10 counter$count = 49412;
	#10 counter$count = 49413;
	#10 counter$count = 49414;
	#10 counter$count = 49415;
	#10 counter$count = 49416;
	#10 counter$count = 49417;
	#10 counter$count = 49418;
	#10 counter$count = 49419;
	#10 counter$count = 49420;
	#10 counter$count = 49421;
	#10 counter$count = 49422;
	#10 counter$count = 49423;
	#10 counter$count = 49424;
	#10 counter$count = 49425;
	#10 counter$count = 49426;
	#10 counter$count = 49427;
	#10 counter$count = 49428;
	#10 counter$count = 49429;
	#10 counter$count = 49430;
	#10 counter$count = 49431;
	#10 counter$count = 49432;
	#10 counter$count = 49433;
	#10 counter$count = 49434;
	#10 counter$count = 49435;
	#10 counter$count = 49436;
	#10 counter$count = 49437;
	#10 counter$count = 49438;
	#10 counter$count = 49439;
	#10 counter$count = 49440;
	#10 counter$count = 49441;
	#10 counter$count = 49442;
	#10 counter$count = 49443;
	#10 counter$count = 49444;
	#10 counter$count = 49445;
	#10 counter$count = 49446;
	#10 counter$count = 49447;
	#10 counter$count = 49448;
	#10 counter$count = 49449;
	#10 counter$count = 49450;
	#10 counter$count = 49451;
	#10 counter$count = 49452;
	#10 counter$count = 49453;
	#10 counter$count = 49454;
	#10 counter$count = 49455;
	#10 counter$count = 49456;
	#10 counter$count = 49457;
	#10 counter$count = 49458;
	#10 counter$count = 49459;
	#10 counter$count = 49460;
	#10 counter$count = 49461;
	#10 counter$count = 49462;
	#10 counter$count = 49463;
	#10 counter$count = 49464;
	#10 counter$count = 49465;
	#10 counter$count = 49466;
	#10 counter$count = 49467;
	#10 counter$count = 49468;
	#10 counter$count = 49469;
	#10 counter$count = 49470;
	#10 counter$count = 49471;
	#10 counter$count = 49472;
	#10 counter$count = 49473;
	#10 counter$count = 49474;
	#10 counter$count = 49475;
	#10 counter$count = 49476;
	#10 counter$count = 49477;
	#10 counter$count = 49478;
	#10 counter$count = 49479;
	#10 counter$count = 49480;
	#10 counter$count = 49481;
	#10 counter$count = 49482;
	#10 counter$count = 49483;
	#10 counter$count = 49484;
	#10 counter$count = 49485;
	#10 counter$count = 49486;
	#10 counter$count = 49487;
	#10 counter$count = 49488;
	#10 counter$count = 49489;
	#10 counter$count = 49490;
	#10 counter$count = 49491;
	#10 counter$count = 49492;
	#10 counter$count = 49493;
	#10 counter$count = 49494;
	#10 counter$count = 49495;
	#10 counter$count = 49496;
	#10 counter$count = 49497;
	#10 counter$count = 49498;
	#10 counter$count = 49499;
	#10 counter$count = 49500;
	#10 counter$count = 49501;
	#10 counter$count = 49502;
	#10 counter$count = 49503;
	#10 counter$count = 49504;
	#10 counter$count = 49505;
	#10 counter$count = 49506;
	#10 counter$count = 49507;
	#10 counter$count = 49508;
	#10 counter$count = 49509;
	#10 counter$count = 49510;
	#10 counter$count = 49511;
	#10 counter$count = 49512;
	#10 counter$count = 49513;
	#10 counter$count = 49514;
	#10 counter$count = 49515;
	#10 counter$count = 49516;
	#10 counter$count = 49517;
	#10 counter$count = 49518;
	#10 counter$count = 49519;
	#10 counter$count = 49520;
	#10 counter$count = 49521;
	#10 counter$count = 49522;
	#10 counter$count = 49523;
	#10 counter$count = 49524;
	#10 counter$count = 49525;
	#10 counter$count = 49526;
	#10 counter$count = 49527;
	#10 counter$count = 49528;
	#10 counter$count = 49529;
	#10 counter$count = 49530;
	#10 counter$count = 49531;
	#10 counter$count = 49532;
	#10 counter$count = 49533;
	#10 counter$count = 49534;
	#10 counter$count = 49535;
	#10 counter$count = 49536;
	#10 counter$count = 49537;
	#10 counter$count = 49538;
	#10 counter$count = 49539;
	#10 counter$count = 49540;
	#10 counter$count = 49541;
	#10 counter$count = 49542;
	#10 counter$count = 49543;
	#10 counter$count = 49544;
	#10 counter$count = 49545;
	#10 counter$count = 49546;
	#10 counter$count = 49547;
	#10 counter$count = 49548;
	#10 counter$count = 49549;
	#10 counter$count = 49550;
	#10 counter$count = 49551;
	#10 counter$count = 49552;
	#10 counter$count = 49553;
	#10 counter$count = 49554;
	#10 counter$count = 49555;
	#10 counter$count = 49556;
	#10 counter$count = 49557;
	#10 counter$count = 49558;
	#10 counter$count = 49559;
	#10 counter$count = 49560;
	#10 counter$count = 49561;
	#10 counter$count = 49562;
	#10 counter$count = 49563;
	#10 counter$count = 49564;
	#10 counter$count = 49565;
	#10 counter$count = 49566;
	#10 counter$count = 49567;
	#10 counter$count = 49568;
	#10 counter$count = 49569;
	#10 counter$count = 49570;
	#10 counter$count = 49571;
	#10 counter$count = 49572;
	#10 counter$count = 49573;
	#10 counter$count = 49574;
	#10 counter$count = 49575;
	#10 counter$count = 49576;
	#10 counter$count = 49577;
	#10 counter$count = 49578;
	#10 counter$count = 49579;
	#10 counter$count = 49580;
	#10 counter$count = 49581;
	#10 counter$count = 49582;
	#10 counter$count = 49583;
	#10 counter$count = 49584;
	#10 counter$count = 49585;
	#10 counter$count = 49586;
	#10 counter$count = 49587;
	#10 counter$count = 49588;
	#10 counter$count = 49589;
	#10 counter$count = 49590;
	#10 counter$count = 49591;
	#10 counter$count = 49592;
	#10 counter$count = 49593;
	#10 counter$count = 49594;
	#10 counter$count = 49595;
	#10 counter$count = 49596;
	#10 counter$count = 49597;
	#10 counter$count = 49598;
	#10 counter$count = 49599;
	#10 counter$count = 49600;
	#10 counter$count = 49601;
	#10 counter$count = 49602;
	#10 counter$count = 49603;
	#10 counter$count = 49604;
	#10 counter$count = 49605;
	#10 counter$count = 49606;
	#10 counter$count = 49607;
	#10 counter$count = 49608;
	#10 counter$count = 49609;
	#10 counter$count = 49610;
	#10 counter$count = 49611;
	#10 counter$count = 49612;
	#10 counter$count = 49613;
	#10 counter$count = 49614;
	#10 counter$count = 49615;
	#10 counter$count = 49616;
	#10 counter$count = 49617;
	#10 counter$count = 49618;
	#10 counter$count = 49619;
	#10 counter$count = 49620;
	#10 counter$count = 49621;
	#10 counter$count = 49622;
	#10 counter$count = 49623;
	#10 counter$count = 49624;
	#10 counter$count = 49625;
	#10 counter$count = 49626;
	#10 counter$count = 49627;
	#10 counter$count = 49628;
	#10 counter$count = 49629;
	#10 counter$count = 49630;
	#10 counter$count = 49631;
	#10 counter$count = 49632;
	#10 counter$count = 49633;
	#10 counter$count = 49634;
	#10 counter$count = 49635;
	#10 counter$count = 49636;
	#10 counter$count = 49637;
	#10 counter$count = 49638;
	#10 counter$count = 49639;
	#10 counter$count = 49640;
	#10 counter$count = 49641;
	#10 counter$count = 49642;
	#10 counter$count = 49643;
	#10 counter$count = 49644;
	#10 counter$count = 49645;
	#10 counter$count = 49646;
	#10 counter$count = 49647;
	#10 counter$count = 49648;
	#10 counter$count = 49649;
	#10 counter$count = 49650;
	#10 counter$count = 49651;
	#10 counter$count = 49652;
	#10 counter$count = 49653;
	#10 counter$count = 49654;
	#10 counter$count = 49655;
	#10 counter$count = 49656;
	#10 counter$count = 49657;
	#10 counter$count = 49658;
	#10 counter$count = 49659;
	#10 counter$count = 49660;
	#10 counter$count = 49661;
	#10 counter$count = 49662;
	#10 counter$count = 49663;
	#10 counter$count = 49664;
	#10 counter$count = 49665;
	#10 counter$count = 49666;
	#10 counter$count = 49667;
	#10 counter$count = 49668;
	#10 counter$count = 49669;
	#10 counter$count = 49670;
	#10 counter$count = 49671;
	#10 counter$count = 49672;
	#10 counter$count = 49673;
	#10 counter$count = 49674;
	#10 counter$count = 49675;
	#10 counter$count = 49676;
	#10 counter$count = 49677;
	#10 counter$count = 49678;
	#10 counter$count = 49679;
	#10 counter$count = 49680;
	#10 counter$count = 49681;
	#10 counter$count = 49682;
	#10 counter$count = 49683;
	#10 counter$count = 49684;
	#10 counter$count = 49685;
	#10 counter$count = 49686;
	#10 counter$count = 49687;
	#10 counter$count = 49688;
	#10 counter$count = 49689;
	#10 counter$count = 49690;
	#10 counter$count = 49691;
	#10 counter$count = 49692;
	#10 counter$count = 49693;
	#10 counter$count = 49694;
	#10 counter$count = 49695;
	#10 counter$count = 49696;
	#10 counter$count = 49697;
	#10 counter$count = 49698;
	#10 counter$count = 49699;
	#10 counter$count = 49700;
	#10 counter$count = 49701;
	#10 counter$count = 49702;
	#10 counter$count = 49703;
	#10 counter$count = 49704;
	#10 counter$count = 49705;
	#10 counter$count = 49706;
	#10 counter$count = 49707;
	#10 counter$count = 49708;
	#10 counter$count = 49709;
	#10 counter$count = 49710;
	#10 counter$count = 49711;
	#10 counter$count = 49712;
	#10 counter$count = 49713;
	#10 counter$count = 49714;
	#10 counter$count = 49715;
	#10 counter$count = 49716;
	#10 counter$count = 49717;
	#10 counter$count = 49718;
	#10 counter$count = 49719;
	#10 counter$count = 49720;
	#10 counter$count = 49721;
	#10 counter$count = 49722;
	#10 counter$count = 49723;
	#10 counter$count = 49724;
	#10 counter$count = 49725;
	#10 counter$count = 49726;
	#10 counter$count = 49727;
	#10 counter$count = 49728;
	#10 counter$count = 49729;
	#10 counter$count = 49730;
	#10 counter$count = 49731;
	#10 counter$count = 49732;
	#10 counter$count = 49733;
	#10 counter$count = 49734;
	#10 counter$count = 49735;
	#10 counter$count = 49736;
	#10 counter$count = 49737;
	#10 counter$count = 49738;
	#10 counter$count = 49739;
	#10 counter$count = 49740;
	#10 counter$count = 49741;
	#10 counter$count = 49742;
	#10 counter$count = 49743;
	#10 counter$count = 49744;
	#10 counter$count = 49745;
	#10 counter$count = 49746;
	#10 counter$count = 49747;
	#10 counter$count = 49748;
	#10 counter$count = 49749;
	#10 counter$count = 49750;
	#10 counter$count = 49751;
	#10 counter$count = 49752;
	#10 counter$count = 49753;
	#10 counter$count = 49754;
	#10 counter$count = 49755;
	#10 counter$count = 49756;
	#10 counter$count = 49757;
	#10 counter$count = 49758;
	#10 counter$count = 49759;
	#10 counter$count = 49760;
	#10 counter$count = 49761;
	#10 counter$count = 49762;
	#10 counter$count = 49763;
	#10 counter$count = 49764;
	#10 counter$count = 49765;
	#10 counter$count = 49766;
	#10 counter$count = 49767;
	#10 counter$count = 49768;
	#10 counter$count = 49769;
	#10 counter$count = 49770;
	#10 counter$count = 49771;
	#10 counter$count = 49772;
	#10 counter$count = 49773;
	#10 counter$count = 49774;
	#10 counter$count = 49775;
	#10 counter$count = 49776;
	#10 counter$count = 49777;
	#10 counter$count = 49778;
	#10 counter$count = 49779;
	#10 counter$count = 49780;
	#10 counter$count = 49781;
	#10 counter$count = 49782;
	#10 counter$count = 49783;
	#10 counter$count = 49784;
	#10 counter$count = 49785;
	#10 counter$count = 49786;
	#10 counter$count = 49787;
	#10 counter$count = 49788;
	#10 counter$count = 49789;
	#10 counter$count = 49790;
	#10 counter$count = 49791;
	#10 counter$count = 49792;
	#10 counter$count = 49793;
	#10 counter$count = 49794;
	#10 counter$count = 49795;
	#10 counter$count = 49796;
	#10 counter$count = 49797;
	#10 counter$count = 49798;
	#10 counter$count = 49799;
	#10 counter$count = 49800;
	#10 counter$count = 49801;
	#10 counter$count = 49802;
	#10 counter$count = 49803;
	#10 counter$count = 49804;
	#10 counter$count = 49805;
	#10 counter$count = 49806;
	#10 counter$count = 49807;
	#10 counter$count = 49808;
	#10 counter$count = 49809;
	#10 counter$count = 49810;
	#10 counter$count = 49811;
	#10 counter$count = 49812;
	#10 counter$count = 49813;
	#10 counter$count = 49814;
	#10 counter$count = 49815;
	#10 counter$count = 49816;
	#10 counter$count = 49817;
	#10 counter$count = 49818;
	#10 counter$count = 49819;
	#10 counter$count = 49820;
	#10 counter$count = 49821;
	#10 counter$count = 49822;
	#10 counter$count = 49823;
	#10 counter$count = 49824;
	#10 counter$count = 49825;
	#10 counter$count = 49826;
	#10 counter$count = 49827;
	#10 counter$count = 49828;
	#10 counter$count = 49829;
	#10 counter$count = 49830;
	#10 counter$count = 49831;
	#10 counter$count = 49832;
	#10 counter$count = 49833;
	#10 counter$count = 49834;
	#10 counter$count = 49835;
	#10 counter$count = 49836;
	#10 counter$count = 49837;
	#10 counter$count = 49838;
	#10 counter$count = 49839;
	#10 counter$count = 49840;
	#10 counter$count = 49841;
	#10 counter$count = 49842;
	#10 counter$count = 49843;
	#10 counter$count = 49844;
	#10 counter$count = 49845;
	#10 counter$count = 49846;
	#10 counter$count = 49847;
	#10 counter$count = 49848;
	#10 counter$count = 49849;
	#10 counter$count = 49850;
	#10 counter$count = 49851;
	#10 counter$count = 49852;
	#10 counter$count = 49853;
	#10 counter$count = 49854;
	#10 counter$count = 49855;
	#10 counter$count = 49856;
	#10 counter$count = 49857;
	#10 counter$count = 49858;
	#10 counter$count = 49859;
	#10 counter$count = 49860;
	#10 counter$count = 49861;
	#10 counter$count = 49862;
	#10 counter$count = 49863;
	#10 counter$count = 49864;
	#10 counter$count = 49865;
	#10 counter$count = 49866;
	#10 counter$count = 49867;
	#10 counter$count = 49868;
	#10 counter$count = 49869;
	#10 counter$count = 49870;
	#10 counter$count = 49871;
	#10 counter$count = 49872;
	#10 counter$count = 49873;
	#10 counter$count = 49874;
	#10 counter$count = 49875;
	#10 counter$count = 49876;
	#10 counter$count = 49877;
	#10 counter$count = 49878;
	#10 counter$count = 49879;
	#10 counter$count = 49880;
	#10 counter$count = 49881;
	#10 counter$count = 49882;
	#10 counter$count = 49883;
	#10 counter$count = 49884;
	#10 counter$count = 49885;
	#10 counter$count = 49886;
	#10 counter$count = 49887;
	#10 counter$count = 49888;
	#10 counter$count = 49889;
	#10 counter$count = 49890;
	#10 counter$count = 49891;
	#10 counter$count = 49892;
	#10 counter$count = 49893;
	#10 counter$count = 49894;
	#10 counter$count = 49895;
	#10 counter$count = 49896;
	#10 counter$count = 49897;
	#10 counter$count = 49898;
	#10 counter$count = 49899;
	#10 counter$count = 49900;
	#10 counter$count = 49901;
	#10 counter$count = 49902;
	#10 counter$count = 49903;
	#10 counter$count = 49904;
	#10 counter$count = 49905;
	#10 counter$count = 49906;
	#10 counter$count = 49907;
	#10 counter$count = 49908;
	#10 counter$count = 49909;
	#10 counter$count = 49910;
	#10 counter$count = 49911;
	#10 counter$count = 49912;
	#10 counter$count = 49913;
	#10 counter$count = 49914;
	#10 counter$count = 49915;
	#10 counter$count = 49916;
	#10 counter$count = 49917;
	#10 counter$count = 49918;
	#10 counter$count = 49919;
	#10 counter$count = 49920;
	#10 counter$count = 49921;
	#10 counter$count = 49922;
	#10 counter$count = 49923;
	#10 counter$count = 49924;
	#10 counter$count = 49925;
	#10 counter$count = 49926;
	#10 counter$count = 49927;
	#10 counter$count = 49928;
	#10 counter$count = 49929;
	#10 counter$count = 49930;
	#10 counter$count = 49931;
	#10 counter$count = 49932;
	#10 counter$count = 49933;
	#10 counter$count = 49934;
	#10 counter$count = 49935;
	#10 counter$count = 49936;
	#10 counter$count = 49937;
	#10 counter$count = 49938;
	#10 counter$count = 49939;
	#10 counter$count = 49940;
	#10 counter$count = 49941;
	#10 counter$count = 49942;
	#10 counter$count = 49943;
	#10 counter$count = 49944;
	#10 counter$count = 49945;
	#10 counter$count = 49946;
	#10 counter$count = 49947;
	#10 counter$count = 49948;
	#10 counter$count = 49949;
	#10 counter$count = 49950;
	#10 counter$count = 49951;
	#10 counter$count = 49952;
	#10 counter$count = 49953;
	#10 counter$count = 49954;
	#10 counter$count = 49955;
	#10 counter$count = 49956;
	#10 counter$count = 49957;
	#10 counter$count = 49958;
	#10 counter$count = 49959;
	#10 counter$count = 49960;
	#10 counter$count = 49961;
	#10 counter$count = 49962;
	#10 counter$count = 49963;
	#10 counter$count = 49964;
	#10 counter$count = 49965;
	#10 counter$count = 49966;
	#10 counter$count = 49967;
	#10 counter$count = 49968;
	#10 counter$count = 49969;
	#10 counter$count = 49970;
	#10 counter$count = 49971;
	#10 counter$count = 49972;
	#10 counter$count = 49973;
	#10 counter$count = 49974;
	#10 counter$count = 49975;
	#10 counter$count = 49976;
	#10 counter$count = 49977;
	#10 counter$count = 49978;
	#10 counter$count = 49979;
	#10 counter$count = 49980;
	#10 counter$count = 49981;
	#10 counter$count = 49982;
	#10 counter$count = 49983;
	#10 counter$count = 49984;
	#10 counter$count = 49985;
	#10 counter$count = 49986;
	#10 counter$count = 49987;
	#10 counter$count = 49988;
	#10 counter$count = 49989;
	#10 counter$count = 49990;
	#10 counter$count = 49991;
	#10 counter$count = 49992;
	#10 counter$count = 49993;
	#10 counter$count = 49994;
	#10 counter$count = 49995;
	#10 counter$count = 49996;
	#10 counter$count = 49997;
	#10 counter$count = 49998;
	#10 counter$count = 49999;
	#10 counter$count = 50000;
	#10 counter$count = 50001;
	#10 counter$count = 50002;
	#10 counter$count = 50003;
	#10 counter$count = 50004;
	#10 counter$count = 50005;
	#10 counter$count = 50006;
	#10 counter$count = 50007;
	#10 counter$count = 50008;
	#10 counter$count = 50009;
	#10 counter$count = 50010;
	#10 counter$count = 50011;
	#10 counter$count = 50012;
	#10 counter$count = 50013;
	#10 counter$count = 50014;
	#10 counter$count = 50015;
	#10 counter$count = 50016;
	#10 counter$count = 50017;
	#10 counter$count = 50018;
	#10 counter$count = 50019;
	#10 counter$count = 50020;
	#10 counter$count = 50021;
	#10 counter$count = 50022;
	#10 counter$count = 50023;
	#10 counter$count = 50024;
	#10 counter$count = 50025;
	#10 counter$count = 50026;
	#10 counter$count = 50027;
	#10 counter$count = 50028;
	#10 counter$count = 50029;
	#10 counter$count = 50030;
	#10 counter$count = 50031;
	#10 counter$count = 50032;
	#10 counter$count = 50033;
	#10 counter$count = 50034;
	#10 counter$count = 50035;
	#10 counter$count = 50036;
	#10 counter$count = 50037;
	#10 counter$count = 50038;
	#10 counter$count = 50039;
	#10 counter$count = 50040;
	#10 counter$count = 50041;
	#10 counter$count = 50042;
	#10 counter$count = 50043;
	#10 counter$count = 50044;
	#10 counter$count = 50045;
	#10 counter$count = 50046;
	#10 counter$count = 50047;
	#10 counter$count = 50048;
	#10 counter$count = 50049;
	#10 counter$count = 50050;
	#10 counter$count = 50051;
	#10 counter$count = 50052;
	#10 counter$count = 50053;
	#10 counter$count = 50054;
	#10 counter$count = 50055;
	#10 counter$count = 50056;
	#10 counter$count = 50057;
	#10 counter$count = 50058;
	#10 counter$count = 50059;
	#10 counter$count = 50060;
	#10 counter$count = 50061;
	#10 counter$count = 50062;
	#10 counter$count = 50063;
	#10 counter$count = 50064;
	#10 counter$count = 50065;
	#10 counter$count = 50066;
	#10 counter$count = 50067;
	#10 counter$count = 50068;
	#10 counter$count = 50069;
	#10 counter$count = 50070;
	#10 counter$count = 50071;
	#10 counter$count = 50072;
	#10 counter$count = 50073;
	#10 counter$count = 50074;
	#10 counter$count = 50075;
	#10 counter$count = 50076;
	#10 counter$count = 50077;
	#10 counter$count = 50078;
	#10 counter$count = 50079;
	#10 counter$count = 50080;
	#10 counter$count = 50081;
	#10 counter$count = 50082;
	#10 counter$count = 50083;
	#10 counter$count = 50084;
	#10 counter$count = 50085;
	#10 counter$count = 50086;
	#10 counter$count = 50087;
	#10 counter$count = 50088;
	#10 counter$count = 50089;
	#10 counter$count = 50090;
	#10 counter$count = 50091;
	#10 counter$count = 50092;
	#10 counter$count = 50093;
	#10 counter$count = 50094;
	#10 counter$count = 50095;
	#10 counter$count = 50096;
	#10 counter$count = 50097;
	#10 counter$count = 50098;
	#10 counter$count = 50099;
	#10 counter$count = 50100;
	#10 counter$count = 50101;
	#10 counter$count = 50102;
	#10 counter$count = 50103;
	#10 counter$count = 50104;
	#10 counter$count = 50105;
	#10 counter$count = 50106;
	#10 counter$count = 50107;
	#10 counter$count = 50108;
	#10 counter$count = 50109;
	#10 counter$count = 50110;
	#10 counter$count = 50111;
	#10 counter$count = 50112;
	#10 counter$count = 50113;
	#10 counter$count = 50114;
	#10 counter$count = 50115;
	#10 counter$count = 50116;
	#10 counter$count = 50117;
	#10 counter$count = 50118;
	#10 counter$count = 50119;
	#10 counter$count = 50120;
	#10 counter$count = 50121;
	#10 counter$count = 50122;
	#10 counter$count = 50123;
	#10 counter$count = 50124;
	#10 counter$count = 50125;
	#10 counter$count = 50126;
	#10 counter$count = 50127;
	#10 counter$count = 50128;
	#10 counter$count = 50129;
	#10 counter$count = 50130;
	#10 counter$count = 50131;
	#10 counter$count = 50132;
	#10 counter$count = 50133;
	#10 counter$count = 50134;
	#10 counter$count = 50135;
	#10 counter$count = 50136;
	#10 counter$count = 50137;
	#10 counter$count = 50138;
	#10 counter$count = 50139;
	#10 counter$count = 50140;
	#10 counter$count = 50141;
	#10 counter$count = 50142;
	#10 counter$count = 50143;
	#10 counter$count = 50144;
	#10 counter$count = 50145;
	#10 counter$count = 50146;
	#10 counter$count = 50147;
	#10 counter$count = 50148;
	#10 counter$count = 50149;
	#10 counter$count = 50150;
	#10 counter$count = 50151;
	#10 counter$count = 50152;
	#10 counter$count = 50153;
	#10 counter$count = 50154;
	#10 counter$count = 50155;
	#10 counter$count = 50156;
	#10 counter$count = 50157;
	#10 counter$count = 50158;
	#10 counter$count = 50159;
	#10 counter$count = 50160;
	#10 counter$count = 50161;
	#10 counter$count = 50162;
	#10 counter$count = 50163;
	#10 counter$count = 50164;
	#10 counter$count = 50165;
	#10 counter$count = 50166;
	#10 counter$count = 50167;
	#10 counter$count = 50168;
	#10 counter$count = 50169;
	#10 counter$count = 50170;
	#10 counter$count = 50171;
	#10 counter$count = 50172;
	#10 counter$count = 50173;
	#10 counter$count = 50174;
	#10 counter$count = 50175;
	#10 counter$count = 50176;
	#10 counter$count = 50177;
	#10 counter$count = 50178;
	#10 counter$count = 50179;
	#10 counter$count = 50180;
	#10 counter$count = 50181;
	#10 counter$count = 50182;
	#10 counter$count = 50183;
	#10 counter$count = 50184;
	#10 counter$count = 50185;
	#10 counter$count = 50186;
	#10 counter$count = 50187;
	#10 counter$count = 50188;
	#10 counter$count = 50189;
	#10 counter$count = 50190;
	#10 counter$count = 50191;
	#10 counter$count = 50192;
	#10 counter$count = 50193;
	#10 counter$count = 50194;
	#10 counter$count = 50195;
	#10 counter$count = 50196;
	#10 counter$count = 50197;
	#10 counter$count = 50198;
	#10 counter$count = 50199;
	#10 counter$count = 50200;
	#10 counter$count = 50201;
	#10 counter$count = 50202;
	#10 counter$count = 50203;
	#10 counter$count = 50204;
	#10 counter$count = 50205;
	#10 counter$count = 50206;
	#10 counter$count = 50207;
	#10 counter$count = 50208;
	#10 counter$count = 50209;
	#10 counter$count = 50210;
	#10 counter$count = 50211;
	#10 counter$count = 50212;
	#10 counter$count = 50213;
	#10 counter$count = 50214;
	#10 counter$count = 50215;
	#10 counter$count = 50216;
	#10 counter$count = 50217;
	#10 counter$count = 50218;
	#10 counter$count = 50219;
	#10 counter$count = 50220;
	#10 counter$count = 50221;
	#10 counter$count = 50222;
	#10 counter$count = 50223;
	#10 counter$count = 50224;
	#10 counter$count = 50225;
	#10 counter$count = 50226;
	#10 counter$count = 50227;
	#10 counter$count = 50228;
	#10 counter$count = 50229;
	#10 counter$count = 50230;
	#10 counter$count = 50231;
	#10 counter$count = 50232;
	#10 counter$count = 50233;
	#10 counter$count = 50234;
	#10 counter$count = 50235;
	#10 counter$count = 50236;
	#10 counter$count = 50237;
	#10 counter$count = 50238;
	#10 counter$count = 50239;
	#10 counter$count = 50240;
	#10 counter$count = 50241;
	#10 counter$count = 50242;
	#10 counter$count = 50243;
	#10 counter$count = 50244;
	#10 counter$count = 50245;
	#10 counter$count = 50246;
	#10 counter$count = 50247;
	#10 counter$count = 50248;
	#10 counter$count = 50249;
	#10 counter$count = 50250;
	#10 counter$count = 50251;
	#10 counter$count = 50252;
	#10 counter$count = 50253;
	#10 counter$count = 50254;
	#10 counter$count = 50255;
	#10 counter$count = 50256;
	#10 counter$count = 50257;
	#10 counter$count = 50258;
	#10 counter$count = 50259;
	#10 counter$count = 50260;
	#10 counter$count = 50261;
	#10 counter$count = 50262;
	#10 counter$count = 50263;
	#10 counter$count = 50264;
	#10 counter$count = 50265;
	#10 counter$count = 50266;
	#10 counter$count = 50267;
	#10 counter$count = 50268;
	#10 counter$count = 50269;
	#10 counter$count = 50270;
	#10 counter$count = 50271;
	#10 counter$count = 50272;
	#10 counter$count = 50273;
	#10 counter$count = 50274;
	#10 counter$count = 50275;
	#10 counter$count = 50276;
	#10 counter$count = 50277;
	#10 counter$count = 50278;
	#10 counter$count = 50279;
	#10 counter$count = 50280;
	#10 counter$count = 50281;
	#10 counter$count = 50282;
	#10 counter$count = 50283;
	#10 counter$count = 50284;
	#10 counter$count = 50285;
	#10 counter$count = 50286;
	#10 counter$count = 50287;
	#10 counter$count = 50288;
	#10 counter$count = 50289;
	#10 counter$count = 50290;
	#10 counter$count = 50291;
	#10 counter$count = 50292;
	#10 counter$count = 50293;
	#10 counter$count = 50294;
	#10 counter$count = 50295;
	#10 counter$count = 50296;
	#10 counter$count = 50297;
	#10 counter$count = 50298;
	#10 counter$count = 50299;
	#10 counter$count = 50300;
	#10 counter$count = 50301;
	#10 counter$count = 50302;
	#10 counter$count = 50303;
	#10 counter$count = 50304;
	#10 counter$count = 50305;
	#10 counter$count = 50306;
	#10 counter$count = 50307;
	#10 counter$count = 50308;
	#10 counter$count = 50309;
	#10 counter$count = 50310;
	#10 counter$count = 50311;
	#10 counter$count = 50312;
	#10 counter$count = 50313;
	#10 counter$count = 50314;
	#10 counter$count = 50315;
	#10 counter$count = 50316;
	#10 counter$count = 50317;
	#10 counter$count = 50318;
	#10 counter$count = 50319;
	#10 counter$count = 50320;
	#10 counter$count = 50321;
	#10 counter$count = 50322;
	#10 counter$count = 50323;
	#10 counter$count = 50324;
	#10 counter$count = 50325;
	#10 counter$count = 50326;
	#10 counter$count = 50327;
	#10 counter$count = 50328;
	#10 counter$count = 50329;
	#10 counter$count = 50330;
	#10 counter$count = 50331;
	#10 counter$count = 50332;
	#10 counter$count = 50333;
	#10 counter$count = 50334;
	#10 counter$count = 50335;
	#10 counter$count = 50336;
	#10 counter$count = 50337;
	#10 counter$count = 50338;
	#10 counter$count = 50339;
	#10 counter$count = 50340;
	#10 counter$count = 50341;
	#10 counter$count = 50342;
	#10 counter$count = 50343;
	#10 counter$count = 50344;
	#10 counter$count = 50345;
	#10 counter$count = 50346;
	#10 counter$count = 50347;
	#10 counter$count = 50348;
	#10 counter$count = 50349;
	#10 counter$count = 50350;
	#10 counter$count = 50351;
	#10 counter$count = 50352;
	#10 counter$count = 50353;
	#10 counter$count = 50354;
	#10 counter$count = 50355;
	#10 counter$count = 50356;
	#10 counter$count = 50357;
	#10 counter$count = 50358;
	#10 counter$count = 50359;
	#10 counter$count = 50360;
	#10 counter$count = 50361;
	#10 counter$count = 50362;
	#10 counter$count = 50363;
	#10 counter$count = 50364;
	#10 counter$count = 50365;
	#10 counter$count = 50366;
	#10 counter$count = 50367;
	#10 counter$count = 50368;
	#10 counter$count = 50369;
	#10 counter$count = 50370;
	#10 counter$count = 50371;
	#10 counter$count = 50372;
	#10 counter$count = 50373;
	#10 counter$count = 50374;
	#10 counter$count = 50375;
	#10 counter$count = 50376;
	#10 counter$count = 50377;
	#10 counter$count = 50378;
	#10 counter$count = 50379;
	#10 counter$count = 50380;
	#10 counter$count = 50381;
	#10 counter$count = 50382;
	#10 counter$count = 50383;
	#10 counter$count = 50384;
	#10 counter$count = 50385;
	#10 counter$count = 50386;
	#10 counter$count = 50387;
	#10 counter$count = 50388;
	#10 counter$count = 50389;
	#10 counter$count = 50390;
	#10 counter$count = 50391;
	#10 counter$count = 50392;
	#10 counter$count = 50393;
	#10 counter$count = 50394;
	#10 counter$count = 50395;
	#10 counter$count = 50396;
	#10 counter$count = 50397;
	#10 counter$count = 50398;
	#10 counter$count = 50399;
	#10 counter$count = 50400;
	#10 counter$count = 50401;
	#10 counter$count = 50402;
	#10 counter$count = 50403;
	#10 counter$count = 50404;
	#10 counter$count = 50405;
	#10 counter$count = 50406;
	#10 counter$count = 50407;
	#10 counter$count = 50408;
	#10 counter$count = 50409;
	#10 counter$count = 50410;
	#10 counter$count = 50411;
	#10 counter$count = 50412;
	#10 counter$count = 50413;
	#10 counter$count = 50414;
	#10 counter$count = 50415;
	#10 counter$count = 50416;
	#10 counter$count = 50417;
	#10 counter$count = 50418;
	#10 counter$count = 50419;
	#10 counter$count = 50420;
	#10 counter$count = 50421;
	#10 counter$count = 50422;
	#10 counter$count = 50423;
	#10 counter$count = 50424;
	#10 counter$count = 50425;
	#10 counter$count = 50426;
	#10 counter$count = 50427;
	#10 counter$count = 50428;
	#10 counter$count = 50429;
	#10 counter$count = 50430;
	#10 counter$count = 50431;
	#10 counter$count = 50432;
	#10 counter$count = 50433;
	#10 counter$count = 50434;
	#10 counter$count = 50435;
	#10 counter$count = 50436;
	#10 counter$count = 50437;
	#10 counter$count = 50438;
	#10 counter$count = 50439;
	#10 counter$count = 50440;
	#10 counter$count = 50441;
	#10 counter$count = 50442;
	#10 counter$count = 50443;
	#10 counter$count = 50444;
	#10 counter$count = 50445;
	#10 counter$count = 50446;
	#10 counter$count = 50447;
	#10 counter$count = 50448;
	#10 counter$count = 50449;
	#10 counter$count = 50450;
	#10 counter$count = 50451;
	#10 counter$count = 50452;
	#10 counter$count = 50453;
	#10 counter$count = 50454;
	#10 counter$count = 50455;
	#10 counter$count = 50456;
	#10 counter$count = 50457;
	#10 counter$count = 50458;
	#10 counter$count = 50459;
	#10 counter$count = 50460;
	#10 counter$count = 50461;
	#10 counter$count = 50462;
	#10 counter$count = 50463;
	#10 counter$count = 50464;
	#10 counter$count = 50465;
	#10 counter$count = 50466;
	#10 counter$count = 50467;
	#10 counter$count = 50468;
	#10 counter$count = 50469;
	#10 counter$count = 50470;
	#10 counter$count = 50471;
	#10 counter$count = 50472;
	#10 counter$count = 50473;
	#10 counter$count = 50474;
	#10 counter$count = 50475;
	#10 counter$count = 50476;
	#10 counter$count = 50477;
	#10 counter$count = 50478;
	#10 counter$count = 50479;
	#10 counter$count = 50480;
	#10 counter$count = 50481;
	#10 counter$count = 50482;
	#10 counter$count = 50483;
	#10 counter$count = 50484;
	#10 counter$count = 50485;
	#10 counter$count = 50486;
	#10 counter$count = 50487;
	#10 counter$count = 50488;
	#10 counter$count = 50489;
	#10 counter$count = 50490;
	#10 counter$count = 50491;
	#10 counter$count = 50492;
	#10 counter$count = 50493;
	#10 counter$count = 50494;
	#10 counter$count = 50495;
	#10 counter$count = 50496;
	#10 counter$count = 50497;
	#10 counter$count = 50498;
	#10 counter$count = 50499;
	#10 counter$count = 50500;
	#10 counter$count = 50501;
	#10 counter$count = 50502;
	#10 counter$count = 50503;
	#10 counter$count = 50504;
	#10 counter$count = 50505;
	#10 counter$count = 50506;
	#10 counter$count = 50507;
	#10 counter$count = 50508;
	#10 counter$count = 50509;
	#10 counter$count = 50510;
	#10 counter$count = 50511;
	#10 counter$count = 50512;
	#10 counter$count = 50513;
	#10 counter$count = 50514;
	#10 counter$count = 50515;
	#10 counter$count = 50516;
	#10 counter$count = 50517;
	#10 counter$count = 50518;
	#10 counter$count = 50519;
	#10 counter$count = 50520;
	#10 counter$count = 50521;
	#10 counter$count = 50522;
	#10 counter$count = 50523;
	#10 counter$count = 50524;
	#10 counter$count = 50525;
	#10 counter$count = 50526;
	#10 counter$count = 50527;
	#10 counter$count = 50528;
	#10 counter$count = 50529;
	#10 counter$count = 50530;
	#10 counter$count = 50531;
	#10 counter$count = 50532;
	#10 counter$count = 50533;
	#10 counter$count = 50534;
	#10 counter$count = 50535;
	#10 counter$count = 50536;
	#10 counter$count = 50537;
	#10 counter$count = 50538;
	#10 counter$count = 50539;
	#10 counter$count = 50540;
	#10 counter$count = 50541;
	#10 counter$count = 50542;
	#10 counter$count = 50543;
	#10 counter$count = 50544;
	#10 counter$count = 50545;
	#10 counter$count = 50546;
	#10 counter$count = 50547;
	#10 counter$count = 50548;
	#10 counter$count = 50549;
	#10 counter$count = 50550;
	#10 counter$count = 50551;
	#10 counter$count = 50552;
	#10 counter$count = 50553;
	#10 counter$count = 50554;
	#10 counter$count = 50555;
	#10 counter$count = 50556;
	#10 counter$count = 50557;
	#10 counter$count = 50558;
	#10 counter$count = 50559;
	#10 counter$count = 50560;
	#10 counter$count = 50561;
	#10 counter$count = 50562;
	#10 counter$count = 50563;
	#10 counter$count = 50564;
	#10 counter$count = 50565;
	#10 counter$count = 50566;
	#10 counter$count = 50567;
	#10 counter$count = 50568;
	#10 counter$count = 50569;
	#10 counter$count = 50570;
	#10 counter$count = 50571;
	#10 counter$count = 50572;
	#10 counter$count = 50573;
	#10 counter$count = 50574;
	#10 counter$count = 50575;
	#10 counter$count = 50576;
	#10 counter$count = 50577;
	#10 counter$count = 50578;
	#10 counter$count = 50579;
	#10 counter$count = 50580;
	#10 counter$count = 50581;
	#10 counter$count = 50582;
	#10 counter$count = 50583;
	#10 counter$count = 50584;
	#10 counter$count = 50585;
	#10 counter$count = 50586;
	#10 counter$count = 50587;
	#10 counter$count = 50588;
	#10 counter$count = 50589;
	#10 counter$count = 50590;
	#10 counter$count = 50591;
	#10 counter$count = 50592;
	#10 counter$count = 50593;
	#10 counter$count = 50594;
	#10 counter$count = 50595;
	#10 counter$count = 50596;
	#10 counter$count = 50597;
	#10 counter$count = 50598;
	#10 counter$count = 50599;
	#10 counter$count = 50600;
	#10 counter$count = 50601;
	#10 counter$count = 50602;
	#10 counter$count = 50603;
	#10 counter$count = 50604;
	#10 counter$count = 50605;
	#10 counter$count = 50606;
	#10 counter$count = 50607;
	#10 counter$count = 50608;
	#10 counter$count = 50609;
	#10 counter$count = 50610;
	#10 counter$count = 50611;
	#10 counter$count = 50612;
	#10 counter$count = 50613;
	#10 counter$count = 50614;
	#10 counter$count = 50615;
	#10 counter$count = 50616;
	#10 counter$count = 50617;
	#10 counter$count = 50618;
	#10 counter$count = 50619;
	#10 counter$count = 50620;
	#10 counter$count = 50621;
	#10 counter$count = 50622;
	#10 counter$count = 50623;
	#10 counter$count = 50624;
	#10 counter$count = 50625;
	#10 counter$count = 50626;
	#10 counter$count = 50627;
	#10 counter$count = 50628;
	#10 counter$count = 50629;
	#10 counter$count = 50630;
	#10 counter$count = 50631;
	#10 counter$count = 50632;
	#10 counter$count = 50633;
	#10 counter$count = 50634;
	#10 counter$count = 50635;
	#10 counter$count = 50636;
	#10 counter$count = 50637;
	#10 counter$count = 50638;
	#10 counter$count = 50639;
	#10 counter$count = 50640;
	#10 counter$count = 50641;
	#10 counter$count = 50642;
	#10 counter$count = 50643;
	#10 counter$count = 50644;
	#10 counter$count = 50645;
	#10 counter$count = 50646;
	#10 counter$count = 50647;
	#10 counter$count = 50648;
	#10 counter$count = 50649;
	#10 counter$count = 50650;
	#10 counter$count = 50651;
	#10 counter$count = 50652;
	#10 counter$count = 50653;
	#10 counter$count = 50654;
	#10 counter$count = 50655;
	#10 counter$count = 50656;
	#10 counter$count = 50657;
	#10 counter$count = 50658;
	#10 counter$count = 50659;
	#10 counter$count = 50660;
	#10 counter$count = 50661;
	#10 counter$count = 50662;
	#10 counter$count = 50663;
	#10 counter$count = 50664;
	#10 counter$count = 50665;
	#10 counter$count = 50666;
	#10 counter$count = 50667;
	#10 counter$count = 50668;
	#10 counter$count = 50669;
	#10 counter$count = 50670;
	#10 counter$count = 50671;
	#10 counter$count = 50672;
	#10 counter$count = 50673;
	#10 counter$count = 50674;
	#10 counter$count = 50675;
	#10 counter$count = 50676;
	#10 counter$count = 50677;
	#10 counter$count = 50678;
	#10 counter$count = 50679;
	#10 counter$count = 50680;
	#10 counter$count = 50681;
	#10 counter$count = 50682;
	#10 counter$count = 50683;
	#10 counter$count = 50684;
	#10 counter$count = 50685;
	#10 counter$count = 50686;
	#10 counter$count = 50687;
	#10 counter$count = 50688;
	#10 counter$count = 50689;
	#10 counter$count = 50690;
	#10 counter$count = 50691;
	#10 counter$count = 50692;
	#10 counter$count = 50693;
	#10 counter$count = 50694;
	#10 counter$count = 50695;
	#10 counter$count = 50696;
	#10 counter$count = 50697;
	#10 counter$count = 50698;
	#10 counter$count = 50699;
	#10 counter$count = 50700;
	#10 counter$count = 50701;
	#10 counter$count = 50702;
	#10 counter$count = 50703;
	#10 counter$count = 50704;
	#10 counter$count = 50705;
	#10 counter$count = 50706;
	#10 counter$count = 50707;
	#10 counter$count = 50708;
	#10 counter$count = 50709;
	#10 counter$count = 50710;
	#10 counter$count = 50711;
	#10 counter$count = 50712;
	#10 counter$count = 50713;
	#10 counter$count = 50714;
	#10 counter$count = 50715;
	#10 counter$count = 50716;
	#10 counter$count = 50717;
	#10 counter$count = 50718;
	#10 counter$count = 50719;
	#10 counter$count = 50720;
	#10 counter$count = 50721;
	#10 counter$count = 50722;
	#10 counter$count = 50723;
	#10 counter$count = 50724;
	#10 counter$count = 50725;
	#10 counter$count = 50726;
	#10 counter$count = 50727;
	#10 counter$count = 50728;
	#10 counter$count = 50729;
	#10 counter$count = 50730;
	#10 counter$count = 50731;
	#10 counter$count = 50732;
	#10 counter$count = 50733;
	#10 counter$count = 50734;
	#10 counter$count = 50735;
	#10 counter$count = 50736;
	#10 counter$count = 50737;
	#10 counter$count = 50738;
	#10 counter$count = 50739;
	#10 counter$count = 50740;
	#10 counter$count = 50741;
	#10 counter$count = 50742;
	#10 counter$count = 50743;
	#10 counter$count = 50744;
	#10 counter$count = 50745;
	#10 counter$count = 50746;
	#10 counter$count = 50747;
	#10 counter$count = 50748;
	#10 counter$count = 50749;
	#10 counter$count = 50750;
	#10 counter$count = 50751;
	#10 counter$count = 50752;
	#10 counter$count = 50753;
	#10 counter$count = 50754;
	#10 counter$count = 50755;
	#10 counter$count = 50756;
	#10 counter$count = 50757;
	#10 counter$count = 50758;
	#10 counter$count = 50759;
	#10 counter$count = 50760;
	#10 counter$count = 50761;
	#10 counter$count = 50762;
	#10 counter$count = 50763;
	#10 counter$count = 50764;
	#10 counter$count = 50765;
	#10 counter$count = 50766;
	#10 counter$count = 50767;
	#10 counter$count = 50768;
	#10 counter$count = 50769;
	#10 counter$count = 50770;
	#10 counter$count = 50771;
	#10 counter$count = 50772;
	#10 counter$count = 50773;
	#10 counter$count = 50774;
	#10 counter$count = 50775;
	#10 counter$count = 50776;
	#10 counter$count = 50777;
	#10 counter$count = 50778;
	#10 counter$count = 50779;
	#10 counter$count = 50780;
	#10 counter$count = 50781;
	#10 counter$count = 50782;
	#10 counter$count = 50783;
	#10 counter$count = 50784;
	#10 counter$count = 50785;
	#10 counter$count = 50786;
	#10 counter$count = 50787;
	#10 counter$count = 50788;
	#10 counter$count = 50789;
	#10 counter$count = 50790;
	#10 counter$count = 50791;
	#10 counter$count = 50792;
	#10 counter$count = 50793;
	#10 counter$count = 50794;
	#10 counter$count = 50795;
	#10 counter$count = 50796;
	#10 counter$count = 50797;
	#10 counter$count = 50798;
	#10 counter$count = 50799;
	#10 counter$count = 50800;
	#10 counter$count = 50801;
	#10 counter$count = 50802;
	#10 counter$count = 50803;
	#10 counter$count = 50804;
	#10 counter$count = 50805;
	#10 counter$count = 50806;
	#10 counter$count = 50807;
	#10 counter$count = 50808;
	#10 counter$count = 50809;
	#10 counter$count = 50810;
	#10 counter$count = 50811;
	#10 counter$count = 50812;
	#10 counter$count = 50813;
	#10 counter$count = 50814;
	#10 counter$count = 50815;
	#10 counter$count = 50816;
	#10 counter$count = 50817;
	#10 counter$count = 50818;
	#10 counter$count = 50819;
	#10 counter$count = 50820;
	#10 counter$count = 50821;
	#10 counter$count = 50822;
	#10 counter$count = 50823;
	#10 counter$count = 50824;
	#10 counter$count = 50825;
	#10 counter$count = 50826;
	#10 counter$count = 50827;
	#10 counter$count = 50828;
	#10 counter$count = 50829;
	#10 counter$count = 50830;
	#10 counter$count = 50831;
	#10 counter$count = 50832;
	#10 counter$count = 50833;
	#10 counter$count = 50834;
	#10 counter$count = 50835;
	#10 counter$count = 50836;
	#10 counter$count = 50837;
	#10 counter$count = 50838;
	#10 counter$count = 50839;
	#10 counter$count = 50840;
	#10 counter$count = 50841;
	#10 counter$count = 50842;
	#10 counter$count = 50843;
	#10 counter$count = 50844;
	#10 counter$count = 50845;
	#10 counter$count = 50846;
	#10 counter$count = 50847;
	#10 counter$count = 50848;
	#10 counter$count = 50849;
	#10 counter$count = 50850;
	#10 counter$count = 50851;
	#10 counter$count = 50852;
	#10 counter$count = 50853;
	#10 counter$count = 50854;
	#10 counter$count = 50855;
	#10 counter$count = 50856;
	#10 counter$count = 50857;
	#10 counter$count = 50858;
	#10 counter$count = 50859;
	#10 counter$count = 50860;
	#10 counter$count = 50861;
	#10 counter$count = 50862;
	#10 counter$count = 50863;
	#10 counter$count = 50864;
	#10 counter$count = 50865;
	#10 counter$count = 50866;
	#10 counter$count = 50867;
	#10 counter$count = 50868;
	#10 counter$count = 50869;
	#10 counter$count = 50870;
	#10 counter$count = 50871;
	#10 counter$count = 50872;
	#10 counter$count = 50873;
	#10 counter$count = 50874;
	#10 counter$count = 50875;
	#10 counter$count = 50876;
	#10 counter$count = 50877;
	#10 counter$count = 50878;
	#10 counter$count = 50879;
	#10 counter$count = 50880;
	#10 counter$count = 50881;
	#10 counter$count = 50882;
	#10 counter$count = 50883;
	#10 counter$count = 50884;
	#10 counter$count = 50885;
	#10 counter$count = 50886;
	#10 counter$count = 50887;
	#10 counter$count = 50888;
	#10 counter$count = 50889;
	#10 counter$count = 50890;
	#10 counter$count = 50891;
	#10 counter$count = 50892;
	#10 counter$count = 50893;
	#10 counter$count = 50894;
	#10 counter$count = 50895;
	#10 counter$count = 50896;
	#10 counter$count = 50897;
	#10 counter$count = 50898;
	#10 counter$count = 50899;
	#10 counter$count = 50900;
	#10 counter$count = 50901;
	#10 counter$count = 50902;
	#10 counter$count = 50903;
	#10 counter$count = 50904;
	#10 counter$count = 50905;
	#10 counter$count = 50906;
	#10 counter$count = 50907;
	#10 counter$count = 50908;
	#10 counter$count = 50909;
	#10 counter$count = 50910;
	#10 counter$count = 50911;
	#10 counter$count = 50912;
	#10 counter$count = 50913;
	#10 counter$count = 50914;
	#10 counter$count = 50915;
	#10 counter$count = 50916;
	#10 counter$count = 50917;
	#10 counter$count = 50918;
	#10 counter$count = 50919;
	#10 counter$count = 50920;
	#10 counter$count = 50921;
	#10 counter$count = 50922;
	#10 counter$count = 50923;
	#10 counter$count = 50924;
	#10 counter$count = 50925;
	#10 counter$count = 50926;
	#10 counter$count = 50927;
	#10 counter$count = 50928;
	#10 counter$count = 50929;
	#10 counter$count = 50930;
	#10 counter$count = 50931;
	#10 counter$count = 50932;
	#10 counter$count = 50933;
	#10 counter$count = 50934;
	#10 counter$count = 50935;
	#10 counter$count = 50936;
	#10 counter$count = 50937;
	#10 counter$count = 50938;
	#10 counter$count = 50939;
	#10 counter$count = 50940;
	#10 counter$count = 50941;
	#10 counter$count = 50942;
	#10 counter$count = 50943;
	#10 counter$count = 50944;
	#10 counter$count = 50945;
	#10 counter$count = 50946;
	#10 counter$count = 50947;
	#10 counter$count = 50948;
	#10 counter$count = 50949;
	#10 counter$count = 50950;
	#10 counter$count = 50951;
	#10 counter$count = 50952;
	#10 counter$count = 50953;
	#10 counter$count = 50954;
	#10 counter$count = 50955;
	#10 counter$count = 50956;
	#10 counter$count = 50957;
	#10 counter$count = 50958;
	#10 counter$count = 50959;
	#10 counter$count = 50960;
	#10 counter$count = 50961;
	#10 counter$count = 50962;
	#10 counter$count = 50963;
	#10 counter$count = 50964;
	#10 counter$count = 50965;
	#10 counter$count = 50966;
	#10 counter$count = 50967;
	#10 counter$count = 50968;
	#10 counter$count = 50969;
	#10 counter$count = 50970;
	#10 counter$count = 50971;
	#10 counter$count = 50972;
	#10 counter$count = 50973;
	#10 counter$count = 50974;
	#10 counter$count = 50975;
	#10 counter$count = 50976;
	#10 counter$count = 50977;
	#10 counter$count = 50978;
	#10 counter$count = 50979;
	#10 counter$count = 50980;
	#10 counter$count = 50981;
	#10 counter$count = 50982;
	#10 counter$count = 50983;
	#10 counter$count = 50984;
	#10 counter$count = 50985;
	#10 counter$count = 50986;
	#10 counter$count = 50987;
	#10 counter$count = 50988;
	#10 counter$count = 50989;
	#10 counter$count = 50990;
	#10 counter$count = 50991;
	#10 counter$count = 50992;
	#10 counter$count = 50993;
	#10 counter$count = 50994;
	#10 counter$count = 50995;
	#10 counter$count = 50996;
	#10 counter$count = 50997;
	#10 counter$count = 50998;
	#10 counter$count = 50999;
	#10 counter$count = 51000;
	#10 counter$count = 51001;
	#10 counter$count = 51002;
	#10 counter$count = 51003;
	#10 counter$count = 51004;
	#10 counter$count = 51005;
	#10 counter$count = 51006;
	#10 counter$count = 51007;
	#10 counter$count = 51008;
	#10 counter$count = 51009;
	#10 counter$count = 51010;
	#10 counter$count = 51011;
	#10 counter$count = 51012;
	#10 counter$count = 51013;
	#10 counter$count = 51014;
	#10 counter$count = 51015;
	#10 counter$count = 51016;
	#10 counter$count = 51017;
	#10 counter$count = 51018;
	#10 counter$count = 51019;
	#10 counter$count = 51020;
	#10 counter$count = 51021;
	#10 counter$count = 51022;
	#10 counter$count = 51023;
	#10 counter$count = 51024;
	#10 counter$count = 51025;
	#10 counter$count = 51026;
	#10 counter$count = 51027;
	#10 counter$count = 51028;
	#10 counter$count = 51029;
	#10 counter$count = 51030;
	#10 counter$count = 51031;
	#10 counter$count = 51032;
	#10 counter$count = 51033;
	#10 counter$count = 51034;
	#10 counter$count = 51035;
	#10 counter$count = 51036;
	#10 counter$count = 51037;
	#10 counter$count = 51038;
	#10 counter$count = 51039;
	#10 counter$count = 51040;
	#10 counter$count = 51041;
	#10 counter$count = 51042;
	#10 counter$count = 51043;
	#10 counter$count = 51044;
	#10 counter$count = 51045;
	#10 counter$count = 51046;
	#10 counter$count = 51047;
	#10 counter$count = 51048;
	#10 counter$count = 51049;
	#10 counter$count = 51050;
	#10 counter$count = 51051;
	#10 counter$count = 51052;
	#10 counter$count = 51053;
	#10 counter$count = 51054;
	#10 counter$count = 51055;
	#10 counter$count = 51056;
	#10 counter$count = 51057;
	#10 counter$count = 51058;
	#10 counter$count = 51059;
	#10 counter$count = 51060;
	#10 counter$count = 51061;
	#10 counter$count = 51062;
	#10 counter$count = 51063;
	#10 counter$count = 51064;
	#10 counter$count = 51065;
	#10 counter$count = 51066;
	#10 counter$count = 51067;
	#10 counter$count = 51068;
	#10 counter$count = 51069;
	#10 counter$count = 51070;
	#10 counter$count = 51071;
	#10 counter$count = 51072;
	#10 counter$count = 51073;
	#10 counter$count = 51074;
	#10 counter$count = 51075;
	#10 counter$count = 51076;
	#10 counter$count = 51077;
	#10 counter$count = 51078;
	#10 counter$count = 51079;
	#10 counter$count = 51080;
	#10 counter$count = 51081;
	#10 counter$count = 51082;
	#10 counter$count = 51083;
	#10 counter$count = 51084;
	#10 counter$count = 51085;
	#10 counter$count = 51086;
	#10 counter$count = 51087;
	#10 counter$count = 51088;
	#10 counter$count = 51089;
	#10 counter$count = 51090;
	#10 counter$count = 51091;
	#10 counter$count = 51092;
	#10 counter$count = 51093;
	#10 counter$count = 51094;
	#10 counter$count = 51095;
	#10 counter$count = 51096;
	#10 counter$count = 51097;
	#10 counter$count = 51098;
	#10 counter$count = 51099;
	#10 counter$count = 51100;
	#10 counter$count = 51101;
	#10 counter$count = 51102;
	#10 counter$count = 51103;
	#10 counter$count = 51104;
	#10 counter$count = 51105;
	#10 counter$count = 51106;
	#10 counter$count = 51107;
	#10 counter$count = 51108;
	#10 counter$count = 51109;
	#10 counter$count = 51110;
	#10 counter$count = 51111;
	#10 counter$count = 51112;
	#10 counter$count = 51113;
	#10 counter$count = 51114;
	#10 counter$count = 51115;
	#10 counter$count = 51116;
	#10 counter$count = 51117;
	#10 counter$count = 51118;
	#10 counter$count = 51119;
	#10 counter$count = 51120;
	#10 counter$count = 51121;
	#10 counter$count = 51122;
	#10 counter$count = 51123;
	#10 counter$count = 51124;
	#10 counter$count = 51125;
	#10 counter$count = 51126;
	#10 counter$count = 51127;
	#10 counter$count = 51128;
	#10 counter$count = 51129;
	#10 counter$count = 51130;
	#10 counter$count = 51131;
	#10 counter$count = 51132;
	#10 counter$count = 51133;
	#10 counter$count = 51134;
	#10 counter$count = 51135;
	#10 counter$count = 51136;
	#10 counter$count = 51137;
	#10 counter$count = 51138;
	#10 counter$count = 51139;
	#10 counter$count = 51140;
	#10 counter$count = 51141;
	#10 counter$count = 51142;
	#10 counter$count = 51143;
	#10 counter$count = 51144;
	#10 counter$count = 51145;
	#10 counter$count = 51146;
	#10 counter$count = 51147;
	#10 counter$count = 51148;
	#10 counter$count = 51149;
	#10 counter$count = 51150;
	#10 counter$count = 51151;
	#10 counter$count = 51152;
	#10 counter$count = 51153;
	#10 counter$count = 51154;
	#10 counter$count = 51155;
	#10 counter$count = 51156;
	#10 counter$count = 51157;
	#10 counter$count = 51158;
	#10 counter$count = 51159;
	#10 counter$count = 51160;
	#10 counter$count = 51161;
	#10 counter$count = 51162;
	#10 counter$count = 51163;
	#10 counter$count = 51164;
	#10 counter$count = 51165;
	#10 counter$count = 51166;
	#10 counter$count = 51167;
	#10 counter$count = 51168;
	#10 counter$count = 51169;
	#10 counter$count = 51170;
	#10 counter$count = 51171;
	#10 counter$count = 51172;
	#10 counter$count = 51173;
	#10 counter$count = 51174;
	#10 counter$count = 51175;
	#10 counter$count = 51176;
	#10 counter$count = 51177;
	#10 counter$count = 51178;
	#10 counter$count = 51179;
	#10 counter$count = 51180;
	#10 counter$count = 51181;
	#10 counter$count = 51182;
	#10 counter$count = 51183;
	#10 counter$count = 51184;
	#10 counter$count = 51185;
	#10 counter$count = 51186;
	#10 counter$count = 51187;
	#10 counter$count = 51188;
	#10 counter$count = 51189;
	#10 counter$count = 51190;
	#10 counter$count = 51191;
	#10 counter$count = 51192;
	#10 counter$count = 51193;
	#10 counter$count = 51194;
	#10 counter$count = 51195;
	#10 counter$count = 51196;
	#10 counter$count = 51197;
	#10 counter$count = 51198;
	#10 counter$count = 51199;
	#10 counter$count = 51200;
	#10 counter$count = 51201;
	#10 counter$count = 51202;
	#10 counter$count = 51203;
	#10 counter$count = 51204;
	#10 counter$count = 51205;
	#10 counter$count = 51206;
	#10 counter$count = 51207;
	#10 counter$count = 51208;
	#10 counter$count = 51209;
	#10 counter$count = 51210;
	#10 counter$count = 51211;
	#10 counter$count = 51212;
	#10 counter$count = 51213;
	#10 counter$count = 51214;
	#10 counter$count = 51215;
	#10 counter$count = 51216;
	#10 counter$count = 51217;
	#10 counter$count = 51218;
	#10 counter$count = 51219;
	#10 counter$count = 51220;
	#10 counter$count = 51221;
	#10 counter$count = 51222;
	#10 counter$count = 51223;
	#10 counter$count = 51224;
	#10 counter$count = 51225;
	#10 counter$count = 51226;
	#10 counter$count = 51227;
	#10 counter$count = 51228;
	#10 counter$count = 51229;
	#10 counter$count = 51230;
	#10 counter$count = 51231;
	#10 counter$count = 51232;
	#10 counter$count = 51233;
	#10 counter$count = 51234;
	#10 counter$count = 51235;
	#10 counter$count = 51236;
	#10 counter$count = 51237;
	#10 counter$count = 51238;
	#10 counter$count = 51239;
	#10 counter$count = 51240;
	#10 counter$count = 51241;
	#10 counter$count = 51242;
	#10 counter$count = 51243;
	#10 counter$count = 51244;
	#10 counter$count = 51245;
	#10 counter$count = 51246;
	#10 counter$count = 51247;
	#10 counter$count = 51248;
	#10 counter$count = 51249;
	#10 counter$count = 51250;
	#10 counter$count = 51251;
	#10 counter$count = 51252;
	#10 counter$count = 51253;
	#10 counter$count = 51254;
	#10 counter$count = 51255;
	#10 counter$count = 51256;
	#10 counter$count = 51257;
	#10 counter$count = 51258;
	#10 counter$count = 51259;
	#10 counter$count = 51260;
	#10 counter$count = 51261;
	#10 counter$count = 51262;
	#10 counter$count = 51263;
	#10 counter$count = 51264;
	#10 counter$count = 51265;
	#10 counter$count = 51266;
	#10 counter$count = 51267;
	#10 counter$count = 51268;
	#10 counter$count = 51269;
	#10 counter$count = 51270;
	#10 counter$count = 51271;
	#10 counter$count = 51272;
	#10 counter$count = 51273;
	#10 counter$count = 51274;
	#10 counter$count = 51275;
	#10 counter$count = 51276;
	#10 counter$count = 51277;
	#10 counter$count = 51278;
	#10 counter$count = 51279;
	#10 counter$count = 51280;
	#10 counter$count = 51281;
	#10 counter$count = 51282;
	#10 counter$count = 51283;
	#10 counter$count = 51284;
	#10 counter$count = 51285;
	#10 counter$count = 51286;
	#10 counter$count = 51287;
	#10 counter$count = 51288;
	#10 counter$count = 51289;
	#10 counter$count = 51290;
	#10 counter$count = 51291;
	#10 counter$count = 51292;
	#10 counter$count = 51293;
	#10 counter$count = 51294;
	#10 counter$count = 51295;
	#10 counter$count = 51296;
	#10 counter$count = 51297;
	#10 counter$count = 51298;
	#10 counter$count = 51299;
	#10 counter$count = 51300;
	#10 counter$count = 51301;
	#10 counter$count = 51302;
	#10 counter$count = 51303;
	#10 counter$count = 51304;
	#10 counter$count = 51305;
	#10 counter$count = 51306;
	#10 counter$count = 51307;
	#10 counter$count = 51308;
	#10 counter$count = 51309;
	#10 counter$count = 51310;
	#10 counter$count = 51311;
	#10 counter$count = 51312;
	#10 counter$count = 51313;
	#10 counter$count = 51314;
	#10 counter$count = 51315;
	#10 counter$count = 51316;
	#10 counter$count = 51317;
	#10 counter$count = 51318;
	#10 counter$count = 51319;
	#10 counter$count = 51320;
	#10 counter$count = 51321;
	#10 counter$count = 51322;
	#10 counter$count = 51323;
	#10 counter$count = 51324;
	#10 counter$count = 51325;
	#10 counter$count = 51326;
	#10 counter$count = 51327;
	#10 counter$count = 51328;
	#10 counter$count = 51329;
	#10 counter$count = 51330;
	#10 counter$count = 51331;
	#10 counter$count = 51332;
	#10 counter$count = 51333;
	#10 counter$count = 51334;
	#10 counter$count = 51335;
	#10 counter$count = 51336;
	#10 counter$count = 51337;
	#10 counter$count = 51338;
	#10 counter$count = 51339;
	#10 counter$count = 51340;
	#10 counter$count = 51341;
	#10 counter$count = 51342;
	#10 counter$count = 51343;
	#10 counter$count = 51344;
	#10 counter$count = 51345;
	#10 counter$count = 51346;
	#10 counter$count = 51347;
	#10 counter$count = 51348;
	#10 counter$count = 51349;
	#10 counter$count = 51350;
	#10 counter$count = 51351;
	#10 counter$count = 51352;
	#10 counter$count = 51353;
	#10 counter$count = 51354;
	#10 counter$count = 51355;
	#10 counter$count = 51356;
	#10 counter$count = 51357;
	#10 counter$count = 51358;
	#10 counter$count = 51359;
	#10 counter$count = 51360;
	#10 counter$count = 51361;
	#10 counter$count = 51362;
	#10 counter$count = 51363;
	#10 counter$count = 51364;
	#10 counter$count = 51365;
	#10 counter$count = 51366;
	#10 counter$count = 51367;
	#10 counter$count = 51368;
	#10 counter$count = 51369;
	#10 counter$count = 51370;
	#10 counter$count = 51371;
	#10 counter$count = 51372;
	#10 counter$count = 51373;
	#10 counter$count = 51374;
	#10 counter$count = 51375;
	#10 counter$count = 51376;
	#10 counter$count = 51377;
	#10 counter$count = 51378;
	#10 counter$count = 51379;
	#10 counter$count = 51380;
	#10 counter$count = 51381;
	#10 counter$count = 51382;
	#10 counter$count = 51383;
	#10 counter$count = 51384;
	#10 counter$count = 51385;
	#10 counter$count = 51386;
	#10 counter$count = 51387;
	#10 counter$count = 51388;
	#10 counter$count = 51389;
	#10 counter$count = 51390;
	#10 counter$count = 51391;
	#10 counter$count = 51392;
	#10 counter$count = 51393;
	#10 counter$count = 51394;
	#10 counter$count = 51395;
	#10 counter$count = 51396;
	#10 counter$count = 51397;
	#10 counter$count = 51398;
	#10 counter$count = 51399;
	#10 counter$count = 51400;
	#10 counter$count = 51401;
	#10 counter$count = 51402;
	#10 counter$count = 51403;
	#10 counter$count = 51404;
	#10 counter$count = 51405;
	#10 counter$count = 51406;
	#10 counter$count = 51407;
	#10 counter$count = 51408;
	#10 counter$count = 51409;
	#10 counter$count = 51410;
	#10 counter$count = 51411;
	#10 counter$count = 51412;
	#10 counter$count = 51413;
	#10 counter$count = 51414;
	#10 counter$count = 51415;
	#10 counter$count = 51416;
	#10 counter$count = 51417;
	#10 counter$count = 51418;
	#10 counter$count = 51419;
	#10 counter$count = 51420;
	#10 counter$count = 51421;
	#10 counter$count = 51422;
	#10 counter$count = 51423;
	#10 counter$count = 51424;
	#10 counter$count = 51425;
	#10 counter$count = 51426;
	#10 counter$count = 51427;
	#10 counter$count = 51428;
	#10 counter$count = 51429;
	#10 counter$count = 51430;
	#10 counter$count = 51431;
	#10 counter$count = 51432;
	#10 counter$count = 51433;
	#10 counter$count = 51434;
	#10 counter$count = 51435;
	#10 counter$count = 51436;
	#10 counter$count = 51437;
	#10 counter$count = 51438;
	#10 counter$count = 51439;
	#10 counter$count = 51440;
	#10 counter$count = 51441;
	#10 counter$count = 51442;
	#10 counter$count = 51443;
	#10 counter$count = 51444;
	#10 counter$count = 51445;
	#10 counter$count = 51446;
	#10 counter$count = 51447;
	#10 counter$count = 51448;
	#10 counter$count = 51449;
	#10 counter$count = 51450;
	#10 counter$count = 51451;
	#10 counter$count = 51452;
	#10 counter$count = 51453;
	#10 counter$count = 51454;
	#10 counter$count = 51455;
	#10 counter$count = 51456;
	#10 counter$count = 51457;
	#10 counter$count = 51458;
	#10 counter$count = 51459;
	#10 counter$count = 51460;
	#10 counter$count = 51461;
	#10 counter$count = 51462;
	#10 counter$count = 51463;
	#10 counter$count = 51464;
	#10 counter$count = 51465;
	#10 counter$count = 51466;
	#10 counter$count = 51467;
	#10 counter$count = 51468;
	#10 counter$count = 51469;
	#10 counter$count = 51470;
	#10 counter$count = 51471;
	#10 counter$count = 51472;
	#10 counter$count = 51473;
	#10 counter$count = 51474;
	#10 counter$count = 51475;
	#10 counter$count = 51476;
	#10 counter$count = 51477;
	#10 counter$count = 51478;
	#10 counter$count = 51479;
	#10 counter$count = 51480;
	#10 counter$count = 51481;
	#10 counter$count = 51482;
	#10 counter$count = 51483;
	#10 counter$count = 51484;
	#10 counter$count = 51485;
	#10 counter$count = 51486;
	#10 counter$count = 51487;
	#10 counter$count = 51488;
	#10 counter$count = 51489;
	#10 counter$count = 51490;
	#10 counter$count = 51491;
	#10 counter$count = 51492;
	#10 counter$count = 51493;
	#10 counter$count = 51494;
	#10 counter$count = 51495;
	#10 counter$count = 51496;
	#10 counter$count = 51497;
	#10 counter$count = 51498;
	#10 counter$count = 51499;
	#10 counter$count = 51500;
	#10 counter$count = 51501;
	#10 counter$count = 51502;
	#10 counter$count = 51503;
	#10 counter$count = 51504;
	#10 counter$count = 51505;
	#10 counter$count = 51506;
	#10 counter$count = 51507;
	#10 counter$count = 51508;
	#10 counter$count = 51509;
	#10 counter$count = 51510;
	#10 counter$count = 51511;
	#10 counter$count = 51512;
	#10 counter$count = 51513;
	#10 counter$count = 51514;
	#10 counter$count = 51515;
	#10 counter$count = 51516;
	#10 counter$count = 51517;
	#10 counter$count = 51518;
	#10 counter$count = 51519;
	#10 counter$count = 51520;
	#10 counter$count = 51521;
	#10 counter$count = 51522;
	#10 counter$count = 51523;
	#10 counter$count = 51524;
	#10 counter$count = 51525;
	#10 counter$count = 51526;
	#10 counter$count = 51527;
	#10 counter$count = 51528;
	#10 counter$count = 51529;
	#10 counter$count = 51530;
	#10 counter$count = 51531;
	#10 counter$count = 51532;
	#10 counter$count = 51533;
	#10 counter$count = 51534;
	#10 counter$count = 51535;
	#10 counter$count = 51536;
	#10 counter$count = 51537;
	#10 counter$count = 51538;
	#10 counter$count = 51539;
	#10 counter$count = 51540;
	#10 counter$count = 51541;
	#10 counter$count = 51542;
	#10 counter$count = 51543;
	#10 counter$count = 51544;
	#10 counter$count = 51545;
	#10 counter$count = 51546;
	#10 counter$count = 51547;
	#10 counter$count = 51548;
	#10 counter$count = 51549;
	#10 counter$count = 51550;
	#10 counter$count = 51551;
	#10 counter$count = 51552;
	#10 counter$count = 51553;
	#10 counter$count = 51554;
	#10 counter$count = 51555;
	#10 counter$count = 51556;
	#10 counter$count = 51557;
	#10 counter$count = 51558;
	#10 counter$count = 51559;
	#10 counter$count = 51560;
	#10 counter$count = 51561;
	#10 counter$count = 51562;
	#10 counter$count = 51563;
	#10 counter$count = 51564;
	#10 counter$count = 51565;
	#10 counter$count = 51566;
	#10 counter$count = 51567;
	#10 counter$count = 51568;
	#10 counter$count = 51569;
	#10 counter$count = 51570;
	#10 counter$count = 51571;
	#10 counter$count = 51572;
	#10 counter$count = 51573;
	#10 counter$count = 51574;
	#10 counter$count = 51575;
	#10 counter$count = 51576;
	#10 counter$count = 51577;
	#10 counter$count = 51578;
	#10 counter$count = 51579;
	#10 counter$count = 51580;
	#10 counter$count = 51581;
	#10 counter$count = 51582;
	#10 counter$count = 51583;
	#10 counter$count = 51584;
	#10 counter$count = 51585;
	#10 counter$count = 51586;
	#10 counter$count = 51587;
	#10 counter$count = 51588;
	#10 counter$count = 51589;
	#10 counter$count = 51590;
	#10 counter$count = 51591;
	#10 counter$count = 51592;
	#10 counter$count = 51593;
	#10 counter$count = 51594;
	#10 counter$count = 51595;
	#10 counter$count = 51596;
	#10 counter$count = 51597;
	#10 counter$count = 51598;
	#10 counter$count = 51599;
	#10 counter$count = 51600;
	#10 counter$count = 51601;
	#10 counter$count = 51602;
	#10 counter$count = 51603;
	#10 counter$count = 51604;
	#10 counter$count = 51605;
	#10 counter$count = 51606;
	#10 counter$count = 51607;
	#10 counter$count = 51608;
	#10 counter$count = 51609;
	#10 counter$count = 51610;
	#10 counter$count = 51611;
	#10 counter$count = 51612;
	#10 counter$count = 51613;
	#10 counter$count = 51614;
	#10 counter$count = 51615;
	#10 counter$count = 51616;
	#10 counter$count = 51617;
	#10 counter$count = 51618;
	#10 counter$count = 51619;
	#10 counter$count = 51620;
	#10 counter$count = 51621;
	#10 counter$count = 51622;
	#10 counter$count = 51623;
	#10 counter$count = 51624;
	#10 counter$count = 51625;
	#10 counter$count = 51626;
	#10 counter$count = 51627;
	#10 counter$count = 51628;
	#10 counter$count = 51629;
	#10 counter$count = 51630;
	#10 counter$count = 51631;
	#10 counter$count = 51632;
	#10 counter$count = 51633;
	#10 counter$count = 51634;
	#10 counter$count = 51635;
	#10 counter$count = 51636;
	#10 counter$count = 51637;
	#10 counter$count = 51638;
	#10 counter$count = 51639;
	#10 counter$count = 51640;
	#10 counter$count = 51641;
	#10 counter$count = 51642;
	#10 counter$count = 51643;
	#10 counter$count = 51644;
	#10 counter$count = 51645;
	#10 counter$count = 51646;
	#10 counter$count = 51647;
	#10 counter$count = 51648;
	#10 counter$count = 51649;
	#10 counter$count = 51650;
	#10 counter$count = 51651;
	#10 counter$count = 51652;
	#10 counter$count = 51653;
	#10 counter$count = 51654;
	#10 counter$count = 51655;
	#10 counter$count = 51656;
	#10 counter$count = 51657;
	#10 counter$count = 51658;
	#10 counter$count = 51659;
	#10 counter$count = 51660;
	#10 counter$count = 51661;
	#10 counter$count = 51662;
	#10 counter$count = 51663;
	#10 counter$count = 51664;
	#10 counter$count = 51665;
	#10 counter$count = 51666;
	#10 counter$count = 51667;
	#10 counter$count = 51668;
	#10 counter$count = 51669;
	#10 counter$count = 51670;
	#10 counter$count = 51671;
	#10 counter$count = 51672;
	#10 counter$count = 51673;
	#10 counter$count = 51674;
	#10 counter$count = 51675;
	#10 counter$count = 51676;
	#10 counter$count = 51677;
	#10 counter$count = 51678;
	#10 counter$count = 51679;
	#10 counter$count = 51680;
	#10 counter$count = 51681;
	#10 counter$count = 51682;
	#10 counter$count = 51683;
	#10 counter$count = 51684;
	#10 counter$count = 51685;
	#10 counter$count = 51686;
	#10 counter$count = 51687;
	#10 counter$count = 51688;
	#10 counter$count = 51689;
	#10 counter$count = 51690;
	#10 counter$count = 51691;
	#10 counter$count = 51692;
	#10 counter$count = 51693;
	#10 counter$count = 51694;
	#10 counter$count = 51695;
	#10 counter$count = 51696;
	#10 counter$count = 51697;
	#10 counter$count = 51698;
	#10 counter$count = 51699;
	#10 counter$count = 51700;
	#10 counter$count = 51701;
	#10 counter$count = 51702;
	#10 counter$count = 51703;
	#10 counter$count = 51704;
	#10 counter$count = 51705;
	#10 counter$count = 51706;
	#10 counter$count = 51707;
	#10 counter$count = 51708;
	#10 counter$count = 51709;
	#10 counter$count = 51710;
	#10 counter$count = 51711;
	#10 counter$count = 51712;
	#10 counter$count = 51713;
	#10 counter$count = 51714;
	#10 counter$count = 51715;
	#10 counter$count = 51716;
	#10 counter$count = 51717;
	#10 counter$count = 51718;
	#10 counter$count = 51719;
	#10 counter$count = 51720;
	#10 counter$count = 51721;
	#10 counter$count = 51722;
	#10 counter$count = 51723;
	#10 counter$count = 51724;
	#10 counter$count = 51725;
	#10 counter$count = 51726;
	#10 counter$count = 51727;
	#10 counter$count = 51728;
	#10 counter$count = 51729;
	#10 counter$count = 51730;
	#10 counter$count = 51731;
	#10 counter$count = 51732;
	#10 counter$count = 51733;
	#10 counter$count = 51734;
	#10 counter$count = 51735;
	#10 counter$count = 51736;
	#10 counter$count = 51737;
	#10 counter$count = 51738;
	#10 counter$count = 51739;
	#10 counter$count = 51740;
	#10 counter$count = 51741;
	#10 counter$count = 51742;
	#10 counter$count = 51743;
	#10 counter$count = 51744;
	#10 counter$count = 51745;
	#10 counter$count = 51746;
	#10 counter$count = 51747;
	#10 counter$count = 51748;
	#10 counter$count = 51749;
	#10 counter$count = 51750;
	#10 counter$count = 51751;
	#10 counter$count = 51752;
	#10 counter$count = 51753;
	#10 counter$count = 51754;
	#10 counter$count = 51755;
	#10 counter$count = 51756;
	#10 counter$count = 51757;
	#10 counter$count = 51758;
	#10 counter$count = 51759;
	#10 counter$count = 51760;
	#10 counter$count = 51761;
	#10 counter$count = 51762;
	#10 counter$count = 51763;
	#10 counter$count = 51764;
	#10 counter$count = 51765;
	#10 counter$count = 51766;
	#10 counter$count = 51767;
	#10 counter$count = 51768;
	#10 counter$count = 51769;
	#10 counter$count = 51770;
	#10 counter$count = 51771;
	#10 counter$count = 51772;
	#10 counter$count = 51773;
	#10 counter$count = 51774;
	#10 counter$count = 51775;
	#10 counter$count = 51776;
	#10 counter$count = 51777;
	#10 counter$count = 51778;
	#10 counter$count = 51779;
	#10 counter$count = 51780;
	#10 counter$count = 51781;
	#10 counter$count = 51782;
	#10 counter$count = 51783;
	#10 counter$count = 51784;
	#10 counter$count = 51785;
	#10 counter$count = 51786;
	#10 counter$count = 51787;
	#10 counter$count = 51788;
	#10 counter$count = 51789;
	#10 counter$count = 51790;
	#10 counter$count = 51791;
	#10 counter$count = 51792;
	#10 counter$count = 51793;
	#10 counter$count = 51794;
	#10 counter$count = 51795;
	#10 counter$count = 51796;
	#10 counter$count = 51797;
	#10 counter$count = 51798;
	#10 counter$count = 51799;
	#10 counter$count = 51800;
	#10 counter$count = 51801;
	#10 counter$count = 51802;
	#10 counter$count = 51803;
	#10 counter$count = 51804;
	#10 counter$count = 51805;
	#10 counter$count = 51806;
	#10 counter$count = 51807;
	#10 counter$count = 51808;
	#10 counter$count = 51809;
	#10 counter$count = 51810;
	#10 counter$count = 51811;
	#10 counter$count = 51812;
	#10 counter$count = 51813;
	#10 counter$count = 51814;
	#10 counter$count = 51815;
	#10 counter$count = 51816;
	#10 counter$count = 51817;
	#10 counter$count = 51818;
	#10 counter$count = 51819;
	#10 counter$count = 51820;
	#10 counter$count = 51821;
	#10 counter$count = 51822;
	#10 counter$count = 51823;
	#10 counter$count = 51824;
	#10 counter$count = 51825;
	#10 counter$count = 51826;
	#10 counter$count = 51827;
	#10 counter$count = 51828;
	#10 counter$count = 51829;
	#10 counter$count = 51830;
	#10 counter$count = 51831;
	#10 counter$count = 51832;
	#10 counter$count = 51833;
	#10 counter$count = 51834;
	#10 counter$count = 51835;
	#10 counter$count = 51836;
	#10 counter$count = 51837;
	#10 counter$count = 51838;
	#10 counter$count = 51839;
	#10 counter$count = 51840;
	#10 counter$count = 51841;
	#10 counter$count = 51842;
	#10 counter$count = 51843;
	#10 counter$count = 51844;
	#10 counter$count = 51845;
	#10 counter$count = 51846;
	#10 counter$count = 51847;
	#10 counter$count = 51848;
	#10 counter$count = 51849;
	#10 counter$count = 51850;
	#10 counter$count = 51851;
	#10 counter$count = 51852;
	#10 counter$count = 51853;
	#10 counter$count = 51854;
	#10 counter$count = 51855;
	#10 counter$count = 51856;
	#10 counter$count = 51857;
	#10 counter$count = 51858;
	#10 counter$count = 51859;
	#10 counter$count = 51860;
	#10 counter$count = 51861;
	#10 counter$count = 51862;
	#10 counter$count = 51863;
	#10 counter$count = 51864;
	#10 counter$count = 51865;
	#10 counter$count = 51866;
	#10 counter$count = 51867;
	#10 counter$count = 51868;
	#10 counter$count = 51869;
	#10 counter$count = 51870;
	#10 counter$count = 51871;
	#10 counter$count = 51872;
	#10 counter$count = 51873;
	#10 counter$count = 51874;
	#10 counter$count = 51875;
	#10 counter$count = 51876;
	#10 counter$count = 51877;
	#10 counter$count = 51878;
	#10 counter$count = 51879;
	#10 counter$count = 51880;
	#10 counter$count = 51881;
	#10 counter$count = 51882;
	#10 counter$count = 51883;
	#10 counter$count = 51884;
	#10 counter$count = 51885;
	#10 counter$count = 51886;
	#10 counter$count = 51887;
	#10 counter$count = 51888;
	#10 counter$count = 51889;
	#10 counter$count = 51890;
	#10 counter$count = 51891;
	#10 counter$count = 51892;
	#10 counter$count = 51893;
	#10 counter$count = 51894;
	#10 counter$count = 51895;
	#10 counter$count = 51896;
	#10 counter$count = 51897;
	#10 counter$count = 51898;
	#10 counter$count = 51899;
	#10 counter$count = 51900;
	#10 counter$count = 51901;
	#10 counter$count = 51902;
	#10 counter$count = 51903;
	#10 counter$count = 51904;
	#10 counter$count = 51905;
	#10 counter$count = 51906;
	#10 counter$count = 51907;
	#10 counter$count = 51908;
	#10 counter$count = 51909;
	#10 counter$count = 51910;
	#10 counter$count = 51911;
	#10 counter$count = 51912;
	#10 counter$count = 51913;
	#10 counter$count = 51914;
	#10 counter$count = 51915;
	#10 counter$count = 51916;
	#10 counter$count = 51917;
	#10 counter$count = 51918;
	#10 counter$count = 51919;
	#10 counter$count = 51920;
	#10 counter$count = 51921;
	#10 counter$count = 51922;
	#10 counter$count = 51923;
	#10 counter$count = 51924;
	#10 counter$count = 51925;
	#10 counter$count = 51926;
	#10 counter$count = 51927;
	#10 counter$count = 51928;
	#10 counter$count = 51929;
	#10 counter$count = 51930;
	#10 counter$count = 51931;
	#10 counter$count = 51932;
	#10 counter$count = 51933;
	#10 counter$count = 51934;
	#10 counter$count = 51935;
	#10 counter$count = 51936;
	#10 counter$count = 51937;
	#10 counter$count = 51938;
	#10 counter$count = 51939;
	#10 counter$count = 51940;
	#10 counter$count = 51941;
	#10 counter$count = 51942;
	#10 counter$count = 51943;
	#10 counter$count = 51944;
	#10 counter$count = 51945;
	#10 counter$count = 51946;
	#10 counter$count = 51947;
	#10 counter$count = 51948;
	#10 counter$count = 51949;
	#10 counter$count = 51950;
	#10 counter$count = 51951;
	#10 counter$count = 51952;
	#10 counter$count = 51953;
	#10 counter$count = 51954;
	#10 counter$count = 51955;
	#10 counter$count = 51956;
	#10 counter$count = 51957;
	#10 counter$count = 51958;
	#10 counter$count = 51959;
	#10 counter$count = 51960;
	#10 counter$count = 51961;
	#10 counter$count = 51962;
	#10 counter$count = 51963;
	#10 counter$count = 51964;
	#10 counter$count = 51965;
	#10 counter$count = 51966;
	#10 counter$count = 51967;
	#10 counter$count = 51968;
	#10 counter$count = 51969;
	#10 counter$count = 51970;
	#10 counter$count = 51971;
	#10 counter$count = 51972;
	#10 counter$count = 51973;
	#10 counter$count = 51974;
	#10 counter$count = 51975;
	#10 counter$count = 51976;
	#10 counter$count = 51977;
	#10 counter$count = 51978;
	#10 counter$count = 51979;
	#10 counter$count = 51980;
	#10 counter$count = 51981;
	#10 counter$count = 51982;
	#10 counter$count = 51983;
	#10 counter$count = 51984;
	#10 counter$count = 51985;
	#10 counter$count = 51986;
	#10 counter$count = 51987;
	#10 counter$count = 51988;
	#10 counter$count = 51989;
	#10 counter$count = 51990;
	#10 counter$count = 51991;
	#10 counter$count = 51992;
	#10 counter$count = 51993;
	#10 counter$count = 51994;
	#10 counter$count = 51995;
	#10 counter$count = 51996;
	#10 counter$count = 51997;
	#10 counter$count = 51998;
	#10 counter$count = 51999;
	#10 counter$count = 52000;
	#10 counter$count = 52001;
	#10 counter$count = 52002;
	#10 counter$count = 52003;
	#10 counter$count = 52004;
	#10 counter$count = 52005;
	#10 counter$count = 52006;
	#10 counter$count = 52007;
	#10 counter$count = 52008;
	#10 counter$count = 52009;
	#10 counter$count = 52010;
	#10 counter$count = 52011;
	#10 counter$count = 52012;
	#10 counter$count = 52013;
	#10 counter$count = 52014;
	#10 counter$count = 52015;
	#10 counter$count = 52016;
	#10 counter$count = 52017;
	#10 counter$count = 52018;
	#10 counter$count = 52019;
	#10 counter$count = 52020;
	#10 counter$count = 52021;
	#10 counter$count = 52022;
	#10 counter$count = 52023;
	#10 counter$count = 52024;
	#10 counter$count = 52025;
	#10 counter$count = 52026;
	#10 counter$count = 52027;
	#10 counter$count = 52028;
	#10 counter$count = 52029;
	#10 counter$count = 52030;
	#10 counter$count = 52031;
	#10 counter$count = 52032;
	#10 counter$count = 52033;
	#10 counter$count = 52034;
	#10 counter$count = 52035;
	#10 counter$count = 52036;
	#10 counter$count = 52037;
	#10 counter$count = 52038;
	#10 counter$count = 52039;
	#10 counter$count = 52040;
	#10 counter$count = 52041;
	#10 counter$count = 52042;
	#10 counter$count = 52043;
	#10 counter$count = 52044;
	#10 counter$count = 52045;
	#10 counter$count = 52046;
	#10 counter$count = 52047;
	#10 counter$count = 52048;
	#10 counter$count = 52049;
	#10 counter$count = 52050;
	#10 counter$count = 52051;
	#10 counter$count = 52052;
	#10 counter$count = 52053;
	#10 counter$count = 52054;
	#10 counter$count = 52055;
	#10 counter$count = 52056;
	#10 counter$count = 52057;
	#10 counter$count = 52058;
	#10 counter$count = 52059;
	#10 counter$count = 52060;
	#10 counter$count = 52061;
	#10 counter$count = 52062;
	#10 counter$count = 52063;
	#10 counter$count = 52064;
	#10 counter$count = 52065;
	#10 counter$count = 52066;
	#10 counter$count = 52067;
	#10 counter$count = 52068;
	#10 counter$count = 52069;
	#10 counter$count = 52070;
	#10 counter$count = 52071;
	#10 counter$count = 52072;
	#10 counter$count = 52073;
	#10 counter$count = 52074;
	#10 counter$count = 52075;
	#10 counter$count = 52076;
	#10 counter$count = 52077;
	#10 counter$count = 52078;
	#10 counter$count = 52079;
	#10 counter$count = 52080;
	#10 counter$count = 52081;
	#10 counter$count = 52082;
	#10 counter$count = 52083;
	#10 counter$count = 52084;
	#10 counter$count = 52085;
	#10 counter$count = 52086;
	#10 counter$count = 52087;
	#10 counter$count = 52088;
	#10 counter$count = 52089;
	#10 counter$count = 52090;
	#10 counter$count = 52091;
	#10 counter$count = 52092;
	#10 counter$count = 52093;
	#10 counter$count = 52094;
	#10 counter$count = 52095;
	#10 counter$count = 52096;
	#10 counter$count = 52097;
	#10 counter$count = 52098;
	#10 counter$count = 52099;
	#10 counter$count = 52100;
	#10 counter$count = 52101;
	#10 counter$count = 52102;
	#10 counter$count = 52103;
	#10 counter$count = 52104;
	#10 counter$count = 52105;
	#10 counter$count = 52106;
	#10 counter$count = 52107;
	#10 counter$count = 52108;
	#10 counter$count = 52109;
	#10 counter$count = 52110;
	#10 counter$count = 52111;
	#10 counter$count = 52112;
	#10 counter$count = 52113;
	#10 counter$count = 52114;
	#10 counter$count = 52115;
	#10 counter$count = 52116;
	#10 counter$count = 52117;
	#10 counter$count = 52118;
	#10 counter$count = 52119;
	#10 counter$count = 52120;
	#10 counter$count = 52121;
	#10 counter$count = 52122;
	#10 counter$count = 52123;
	#10 counter$count = 52124;
	#10 counter$count = 52125;
	#10 counter$count = 52126;
	#10 counter$count = 52127;
	#10 counter$count = 52128;
	#10 counter$count = 52129;
	#10 counter$count = 52130;
	#10 counter$count = 52131;
	#10 counter$count = 52132;
	#10 counter$count = 52133;
	#10 counter$count = 52134;
	#10 counter$count = 52135;
	#10 counter$count = 52136;
	#10 counter$count = 52137;
	#10 counter$count = 52138;
	#10 counter$count = 52139;
	#10 counter$count = 52140;
	#10 counter$count = 52141;
	#10 counter$count = 52142;
	#10 counter$count = 52143;
	#10 counter$count = 52144;
	#10 counter$count = 52145;
	#10 counter$count = 52146;
	#10 counter$count = 52147;
	#10 counter$count = 52148;
	#10 counter$count = 52149;
	#10 counter$count = 52150;
	#10 counter$count = 52151;
	#10 counter$count = 52152;
	#10 counter$count = 52153;
	#10 counter$count = 52154;
	#10 counter$count = 52155;
	#10 counter$count = 52156;
	#10 counter$count = 52157;
	#10 counter$count = 52158;
	#10 counter$count = 52159;
	#10 counter$count = 52160;
	#10 counter$count = 52161;
	#10 counter$count = 52162;
	#10 counter$count = 52163;
	#10 counter$count = 52164;
	#10 counter$count = 52165;
	#10 counter$count = 52166;
	#10 counter$count = 52167;
	#10 counter$count = 52168;
	#10 counter$count = 52169;
	#10 counter$count = 52170;
	#10 counter$count = 52171;
	#10 counter$count = 52172;
	#10 counter$count = 52173;
	#10 counter$count = 52174;
	#10 counter$count = 52175;
	#10 counter$count = 52176;
	#10 counter$count = 52177;
	#10 counter$count = 52178;
	#10 counter$count = 52179;
	#10 counter$count = 52180;
	#10 counter$count = 52181;
	#10 counter$count = 52182;
	#10 counter$count = 52183;
	#10 counter$count = 52184;
	#10 counter$count = 52185;
	#10 counter$count = 52186;
	#10 counter$count = 52187;
	#10 counter$count = 52188;
	#10 counter$count = 52189;
	#10 counter$count = 52190;
	#10 counter$count = 52191;
	#10 counter$count = 52192;
	#10 counter$count = 52193;
	#10 counter$count = 52194;
	#10 counter$count = 52195;
	#10 counter$count = 52196;
	#10 counter$count = 52197;
	#10 counter$count = 52198;
	#10 counter$count = 52199;
	#10 counter$count = 52200;
	#10 counter$count = 52201;
	#10 counter$count = 52202;
	#10 counter$count = 52203;
	#10 counter$count = 52204;
	#10 counter$count = 52205;
	#10 counter$count = 52206;
	#10 counter$count = 52207;
	#10 counter$count = 52208;
	#10 counter$count = 52209;
	#10 counter$count = 52210;
	#10 counter$count = 52211;
	#10 counter$count = 52212;
	#10 counter$count = 52213;
	#10 counter$count = 52214;
	#10 counter$count = 52215;
	#10 counter$count = 52216;
	#10 counter$count = 52217;
	#10 counter$count = 52218;
	#10 counter$count = 52219;
	#10 counter$count = 52220;
	#10 counter$count = 52221;
	#10 counter$count = 52222;
	#10 counter$count = 52223;
	#10 counter$count = 52224;
	#10 counter$count = 52225;
	#10 counter$count = 52226;
	#10 counter$count = 52227;
	#10 counter$count = 52228;
	#10 counter$count = 52229;
	#10 counter$count = 52230;
	#10 counter$count = 52231;
	#10 counter$count = 52232;
	#10 counter$count = 52233;
	#10 counter$count = 52234;
	#10 counter$count = 52235;
	#10 counter$count = 52236;
	#10 counter$count = 52237;
	#10 counter$count = 52238;
	#10 counter$count = 52239;
	#10 counter$count = 52240;
	#10 counter$count = 52241;
	#10 counter$count = 52242;
	#10 counter$count = 52243;
	#10 counter$count = 52244;
	#10 counter$count = 52245;
	#10 counter$count = 52246;
	#10 counter$count = 52247;
	#10 counter$count = 52248;
	#10 counter$count = 52249;
	#10 counter$count = 52250;
	#10 counter$count = 52251;
	#10 counter$count = 52252;
	#10 counter$count = 52253;
	#10 counter$count = 52254;
	#10 counter$count = 52255;
	#10 counter$count = 52256;
	#10 counter$count = 52257;
	#10 counter$count = 52258;
	#10 counter$count = 52259;
	#10 counter$count = 52260;
	#10 counter$count = 52261;
	#10 counter$count = 52262;
	#10 counter$count = 52263;
	#10 counter$count = 52264;
	#10 counter$count = 52265;
	#10 counter$count = 52266;
	#10 counter$count = 52267;
	#10 counter$count = 52268;
	#10 counter$count = 52269;
	#10 counter$count = 52270;
	#10 counter$count = 52271;
	#10 counter$count = 52272;
	#10 counter$count = 52273;
	#10 counter$count = 52274;
	#10 counter$count = 52275;
	#10 counter$count = 52276;
	#10 counter$count = 52277;
	#10 counter$count = 52278;
	#10 counter$count = 52279;
	#10 counter$count = 52280;
	#10 counter$count = 52281;
	#10 counter$count = 52282;
	#10 counter$count = 52283;
	#10 counter$count = 52284;
	#10 counter$count = 52285;
	#10 counter$count = 52286;
	#10 counter$count = 52287;
	#10 counter$count = 52288;
	#10 counter$count = 52289;
	#10 counter$count = 52290;
	#10 counter$count = 52291;
	#10 counter$count = 52292;
	#10 counter$count = 52293;
	#10 counter$count = 52294;
	#10 counter$count = 52295;
	#10 counter$count = 52296;
	#10 counter$count = 52297;
	#10 counter$count = 52298;
	#10 counter$count = 52299;
	#10 counter$count = 52300;
	#10 counter$count = 52301;
	#10 counter$count = 52302;
	#10 counter$count = 52303;
	#10 counter$count = 52304;
	#10 counter$count = 52305;
	#10 counter$count = 52306;
	#10 counter$count = 52307;
	#10 counter$count = 52308;
	#10 counter$count = 52309;
	#10 counter$count = 52310;
	#10 counter$count = 52311;
	#10 counter$count = 52312;
	#10 counter$count = 52313;
	#10 counter$count = 52314;
	#10 counter$count = 52315;
	#10 counter$count = 52316;
	#10 counter$count = 52317;
	#10 counter$count = 52318;
	#10 counter$count = 52319;
	#10 counter$count = 52320;
	#10 counter$count = 52321;
	#10 counter$count = 52322;
	#10 counter$count = 52323;
	#10 counter$count = 52324;
	#10 counter$count = 52325;
	#10 counter$count = 52326;
	#10 counter$count = 52327;
	#10 counter$count = 52328;
	#10 counter$count = 52329;
	#10 counter$count = 52330;
	#10 counter$count = 52331;
	#10 counter$count = 52332;
	#10 counter$count = 52333;
	#10 counter$count = 52334;
	#10 counter$count = 52335;
	#10 counter$count = 52336;
	#10 counter$count = 52337;
	#10 counter$count = 52338;
	#10 counter$count = 52339;
	#10 counter$count = 52340;
	#10 counter$count = 52341;
	#10 counter$count = 52342;
	#10 counter$count = 52343;
	#10 counter$count = 52344;
	#10 counter$count = 52345;
	#10 counter$count = 52346;
	#10 counter$count = 52347;
	#10 counter$count = 52348;
	#10 counter$count = 52349;
	#10 counter$count = 52350;
	#10 counter$count = 52351;
	#10 counter$count = 52352;
	#10 counter$count = 52353;
	#10 counter$count = 52354;
	#10 counter$count = 52355;
	#10 counter$count = 52356;
	#10 counter$count = 52357;
	#10 counter$count = 52358;
	#10 counter$count = 52359;
	#10 counter$count = 52360;
	#10 counter$count = 52361;
	#10 counter$count = 52362;
	#10 counter$count = 52363;
	#10 counter$count = 52364;
	#10 counter$count = 52365;
	#10 counter$count = 52366;
	#10 counter$count = 52367;
	#10 counter$count = 52368;
	#10 counter$count = 52369;
	#10 counter$count = 52370;
	#10 counter$count = 52371;
	#10 counter$count = 52372;
	#10 counter$count = 52373;
	#10 counter$count = 52374;
	#10 counter$count = 52375;
	#10 counter$count = 52376;
	#10 counter$count = 52377;
	#10 counter$count = 52378;
	#10 counter$count = 52379;
	#10 counter$count = 52380;
	#10 counter$count = 52381;
	#10 counter$count = 52382;
	#10 counter$count = 52383;
	#10 counter$count = 52384;
	#10 counter$count = 52385;
	#10 counter$count = 52386;
	#10 counter$count = 52387;
	#10 counter$count = 52388;
	#10 counter$count = 52389;
	#10 counter$count = 52390;
	#10 counter$count = 52391;
	#10 counter$count = 52392;
	#10 counter$count = 52393;
	#10 counter$count = 52394;
	#10 counter$count = 52395;
	#10 counter$count = 52396;
	#10 counter$count = 52397;
	#10 counter$count = 52398;
	#10 counter$count = 52399;
	#10 counter$count = 52400;
	#10 counter$count = 52401;
	#10 counter$count = 52402;
	#10 counter$count = 52403;
	#10 counter$count = 52404;
	#10 counter$count = 52405;
	#10 counter$count = 52406;
	#10 counter$count = 52407;
	#10 counter$count = 52408;
	#10 counter$count = 52409;
	#10 counter$count = 52410;
	#10 counter$count = 52411;
	#10 counter$count = 52412;
	#10 counter$count = 52413;
	#10 counter$count = 52414;
	#10 counter$count = 52415;
	#10 counter$count = 52416;
	#10 counter$count = 52417;
	#10 counter$count = 52418;
	#10 counter$count = 52419;
	#10 counter$count = 52420;
	#10 counter$count = 52421;
	#10 counter$count = 52422;
	#10 counter$count = 52423;
	#10 counter$count = 52424;
	#10 counter$count = 52425;
	#10 counter$count = 52426;
	#10 counter$count = 52427;
	#10 counter$count = 52428;
	#10 counter$count = 52429;
	#10 counter$count = 52430;
	#10 counter$count = 52431;
	#10 counter$count = 52432;
	#10 counter$count = 52433;
	#10 counter$count = 52434;
	#10 counter$count = 52435;
	#10 counter$count = 52436;
	#10 counter$count = 52437;
	#10 counter$count = 52438;
	#10 counter$count = 52439;
	#10 counter$count = 52440;
	#10 counter$count = 52441;
	#10 counter$count = 52442;
	#10 counter$count = 52443;
	#10 counter$count = 52444;
	#10 counter$count = 52445;
	#10 counter$count = 52446;
	#10 counter$count = 52447;
	#10 counter$count = 52448;
	#10 counter$count = 52449;
	#10 counter$count = 52450;
	#10 counter$count = 52451;
	#10 counter$count = 52452;
	#10 counter$count = 52453;
	#10 counter$count = 52454;
	#10 counter$count = 52455;
	#10 counter$count = 52456;
	#10 counter$count = 52457;
	#10 counter$count = 52458;
	#10 counter$count = 52459;
	#10 counter$count = 52460;
	#10 counter$count = 52461;
	#10 counter$count = 52462;
	#10 counter$count = 52463;
	#10 counter$count = 52464;
	#10 counter$count = 52465;
	#10 counter$count = 52466;
	#10 counter$count = 52467;
	#10 counter$count = 52468;
	#10 counter$count = 52469;
	#10 counter$count = 52470;
	#10 counter$count = 52471;
	#10 counter$count = 52472;
	#10 counter$count = 52473;
	#10 counter$count = 52474;
	#10 counter$count = 52475;
	#10 counter$count = 52476;
	#10 counter$count = 52477;
	#10 counter$count = 52478;
	#10 counter$count = 52479;
	#10 counter$count = 52480;
	#10 counter$count = 52481;
	#10 counter$count = 52482;
	#10 counter$count = 52483;
	#10 counter$count = 52484;
	#10 counter$count = 52485;
	#10 counter$count = 52486;
	#10 counter$count = 52487;
	#10 counter$count = 52488;
	#10 counter$count = 52489;
	#10 counter$count = 52490;
	#10 counter$count = 52491;
	#10 counter$count = 52492;
	#10 counter$count = 52493;
	#10 counter$count = 52494;
	#10 counter$count = 52495;
	#10 counter$count = 52496;
	#10 counter$count = 52497;
	#10 counter$count = 52498;
	#10 counter$count = 52499;
	#10 counter$count = 52500;
	#10 counter$count = 52501;
	#10 counter$count = 52502;
	#10 counter$count = 52503;
	#10 counter$count = 52504;
	#10 counter$count = 52505;
	#10 counter$count = 52506;
	#10 counter$count = 52507;
	#10 counter$count = 52508;
	#10 counter$count = 52509;
	#10 counter$count = 52510;
	#10 counter$count = 52511;
	#10 counter$count = 52512;
	#10 counter$count = 52513;
	#10 counter$count = 52514;
	#10 counter$count = 52515;
	#10 counter$count = 52516;
	#10 counter$count = 52517;
	#10 counter$count = 52518;
	#10 counter$count = 52519;
	#10 counter$count = 52520;
	#10 counter$count = 52521;
	#10 counter$count = 52522;
	#10 counter$count = 52523;
	#10 counter$count = 52524;
	#10 counter$count = 52525;
	#10 counter$count = 52526;
	#10 counter$count = 52527;
	#10 counter$count = 52528;
	#10 counter$count = 52529;
	#10 counter$count = 52530;
	#10 counter$count = 52531;
	#10 counter$count = 52532;
	#10 counter$count = 52533;
	#10 counter$count = 52534;
	#10 counter$count = 52535;
	#10 counter$count = 52536;
	#10 counter$count = 52537;
	#10 counter$count = 52538;
	#10 counter$count = 52539;
	#10 counter$count = 52540;
	#10 counter$count = 52541;
	#10 counter$count = 52542;
	#10 counter$count = 52543;
	#10 counter$count = 52544;
	#10 counter$count = 52545;
	#10 counter$count = 52546;
	#10 counter$count = 52547;
	#10 counter$count = 52548;
	#10 counter$count = 52549;
	#10 counter$count = 52550;
	#10 counter$count = 52551;
	#10 counter$count = 52552;
	#10 counter$count = 52553;
	#10 counter$count = 52554;
	#10 counter$count = 52555;
	#10 counter$count = 52556;
	#10 counter$count = 52557;
	#10 counter$count = 52558;
	#10 counter$count = 52559;
	#10 counter$count = 52560;
	#10 counter$count = 52561;
	#10 counter$count = 52562;
	#10 counter$count = 52563;
	#10 counter$count = 52564;
	#10 counter$count = 52565;
	#10 counter$count = 52566;
	#10 counter$count = 52567;
	#10 counter$count = 52568;
	#10 counter$count = 52569;
	#10 counter$count = 52570;
	#10 counter$count = 52571;
	#10 counter$count = 52572;
	#10 counter$count = 52573;
	#10 counter$count = 52574;
	#10 counter$count = 52575;
	#10 counter$count = 52576;
	#10 counter$count = 52577;
	#10 counter$count = 52578;
	#10 counter$count = 52579;
	#10 counter$count = 52580;
	#10 counter$count = 52581;
	#10 counter$count = 52582;
	#10 counter$count = 52583;
	#10 counter$count = 52584;
	#10 counter$count = 52585;
	#10 counter$count = 52586;
	#10 counter$count = 52587;
	#10 counter$count = 52588;
	#10 counter$count = 52589;
	#10 counter$count = 52590;
	#10 counter$count = 52591;
	#10 counter$count = 52592;
	#10 counter$count = 52593;
	#10 counter$count = 52594;
	#10 counter$count = 52595;
	#10 counter$count = 52596;
	#10 counter$count = 52597;
	#10 counter$count = 52598;
	#10 counter$count = 52599;
	#10 counter$count = 52600;
	#10 counter$count = 52601;
	#10 counter$count = 52602;
	#10 counter$count = 52603;
	#10 counter$count = 52604;
	#10 counter$count = 52605;
	#10 counter$count = 52606;
	#10 counter$count = 52607;
	#10 counter$count = 52608;
	#10 counter$count = 52609;
	#10 counter$count = 52610;
	#10 counter$count = 52611;
	#10 counter$count = 52612;
	#10 counter$count = 52613;
	#10 counter$count = 52614;
	#10 counter$count = 52615;
	#10 counter$count = 52616;
	#10 counter$count = 52617;
	#10 counter$count = 52618;
	#10 counter$count = 52619;
	#10 counter$count = 52620;
	#10 counter$count = 52621;
	#10 counter$count = 52622;
	#10 counter$count = 52623;
	#10 counter$count = 52624;
	#10 counter$count = 52625;
	#10 counter$count = 52626;
	#10 counter$count = 52627;
	#10 counter$count = 52628;
	#10 counter$count = 52629;
	#10 counter$count = 52630;
	#10 counter$count = 52631;
	#10 counter$count = 52632;
	#10 counter$count = 52633;
	#10 counter$count = 52634;
	#10 counter$count = 52635;
	#10 counter$count = 52636;
	#10 counter$count = 52637;
	#10 counter$count = 52638;
	#10 counter$count = 52639;
	#10 counter$count = 52640;
	#10 counter$count = 52641;
	#10 counter$count = 52642;
	#10 counter$count = 52643;
	#10 counter$count = 52644;
	#10 counter$count = 52645;
	#10 counter$count = 52646;
	#10 counter$count = 52647;
	#10 counter$count = 52648;
	#10 counter$count = 52649;
	#10 counter$count = 52650;
	#10 counter$count = 52651;
	#10 counter$count = 52652;
	#10 counter$count = 52653;
	#10 counter$count = 52654;
	#10 counter$count = 52655;
	#10 counter$count = 52656;
	#10 counter$count = 52657;
	#10 counter$count = 52658;
	#10 counter$count = 52659;
	#10 counter$count = 52660;
	#10 counter$count = 52661;
	#10 counter$count = 52662;
	#10 counter$count = 52663;
	#10 counter$count = 52664;
	#10 counter$count = 52665;
	#10 counter$count = 52666;
	#10 counter$count = 52667;
	#10 counter$count = 52668;
	#10 counter$count = 52669;
	#10 counter$count = 52670;
	#10 counter$count = 52671;
	#10 counter$count = 52672;
	#10 counter$count = 52673;
	#10 counter$count = 52674;
	#10 counter$count = 52675;
	#10 counter$count = 52676;
	#10 counter$count = 52677;
	#10 counter$count = 52678;
	#10 counter$count = 52679;
	#10 counter$count = 52680;
	#10 counter$count = 52681;
	#10 counter$count = 52682;
	#10 counter$count = 52683;
	#10 counter$count = 52684;
	#10 counter$count = 52685;
	#10 counter$count = 52686;
	#10 counter$count = 52687;
	#10 counter$count = 52688;
	#10 counter$count = 52689;
	#10 counter$count = 52690;
	#10 counter$count = 52691;
	#10 counter$count = 52692;
	#10 counter$count = 52693;
	#10 counter$count = 52694;
	#10 counter$count = 52695;
	#10 counter$count = 52696;
	#10 counter$count = 52697;
	#10 counter$count = 52698;
	#10 counter$count = 52699;
	#10 counter$count = 52700;
	#10 counter$count = 52701;
	#10 counter$count = 52702;
	#10 counter$count = 52703;
	#10 counter$count = 52704;
	#10 counter$count = 52705;
	#10 counter$count = 52706;
	#10 counter$count = 52707;
	#10 counter$count = 52708;
	#10 counter$count = 52709;
	#10 counter$count = 52710;
	#10 counter$count = 52711;
	#10 counter$count = 52712;
	#10 counter$count = 52713;
	#10 counter$count = 52714;
	#10 counter$count = 52715;
	#10 counter$count = 52716;
	#10 counter$count = 52717;
	#10 counter$count = 52718;
	#10 counter$count = 52719;
	#10 counter$count = 52720;
	#10 counter$count = 52721;
	#10 counter$count = 52722;
	#10 counter$count = 52723;
	#10 counter$count = 52724;
	#10 counter$count = 52725;
	#10 counter$count = 52726;
	#10 counter$count = 52727;
	#10 counter$count = 52728;
	#10 counter$count = 52729;
	#10 counter$count = 52730;
	#10 counter$count = 52731;
	#10 counter$count = 52732;
	#10 counter$count = 52733;
	#10 counter$count = 52734;
	#10 counter$count = 52735;
	#10 counter$count = 52736;
	#10 counter$count = 52737;
	#10 counter$count = 52738;
	#10 counter$count = 52739;
	#10 counter$count = 52740;
	#10 counter$count = 52741;
	#10 counter$count = 52742;
	#10 counter$count = 52743;
	#10 counter$count = 52744;
	#10 counter$count = 52745;
	#10 counter$count = 52746;
	#10 counter$count = 52747;
	#10 counter$count = 52748;
	#10 counter$count = 52749;
	#10 counter$count = 52750;
	#10 counter$count = 52751;
	#10 counter$count = 52752;
	#10 counter$count = 52753;
	#10 counter$count = 52754;
	#10 counter$count = 52755;
	#10 counter$count = 52756;
	#10 counter$count = 52757;
	#10 counter$count = 52758;
	#10 counter$count = 52759;
	#10 counter$count = 52760;
	#10 counter$count = 52761;
	#10 counter$count = 52762;
	#10 counter$count = 52763;
	#10 counter$count = 52764;
	#10 counter$count = 52765;
	#10 counter$count = 52766;
	#10 counter$count = 52767;
	#10 counter$count = 52768;
	#10 counter$count = 52769;
	#10 counter$count = 52770;
	#10 counter$count = 52771;
	#10 counter$count = 52772;
	#10 counter$count = 52773;
	#10 counter$count = 52774;
	#10 counter$count = 52775;
	#10 counter$count = 52776;
	#10 counter$count = 52777;
	#10 counter$count = 52778;
	#10 counter$count = 52779;
	#10 counter$count = 52780;
	#10 counter$count = 52781;
	#10 counter$count = 52782;
	#10 counter$count = 52783;
	#10 counter$count = 52784;
	#10 counter$count = 52785;
	#10 counter$count = 52786;
	#10 counter$count = 52787;
	#10 counter$count = 52788;
	#10 counter$count = 52789;
	#10 counter$count = 52790;
	#10 counter$count = 52791;
	#10 counter$count = 52792;
	#10 counter$count = 52793;
	#10 counter$count = 52794;
	#10 counter$count = 52795;
	#10 counter$count = 52796;
	#10 counter$count = 52797;
	#10 counter$count = 52798;
	#10 counter$count = 52799;
	#10 counter$count = 52800;
	#10 counter$count = 52801;
	#10 counter$count = 52802;
	#10 counter$count = 52803;
	#10 counter$count = 52804;
	#10 counter$count = 52805;
	#10 counter$count = 52806;
	#10 counter$count = 52807;
	#10 counter$count = 52808;
	#10 counter$count = 52809;
	#10 counter$count = 52810;
	#10 counter$count = 52811;
	#10 counter$count = 52812;
	#10 counter$count = 52813;
	#10 counter$count = 52814;
	#10 counter$count = 52815;
	#10 counter$count = 52816;
	#10 counter$count = 52817;
	#10 counter$count = 52818;
	#10 counter$count = 52819;
	#10 counter$count = 52820;
	#10 counter$count = 52821;
	#10 counter$count = 52822;
	#10 counter$count = 52823;
	#10 counter$count = 52824;
	#10 counter$count = 52825;
	#10 counter$count = 52826;
	#10 counter$count = 52827;
	#10 counter$count = 52828;
	#10 counter$count = 52829;
	#10 counter$count = 52830;
	#10 counter$count = 52831;
	#10 counter$count = 52832;
	#10 counter$count = 52833;
	#10 counter$count = 52834;
	#10 counter$count = 52835;
	#10 counter$count = 52836;
	#10 counter$count = 52837;
	#10 counter$count = 52838;
	#10 counter$count = 52839;
	#10 counter$count = 52840;
	#10 counter$count = 52841;
	#10 counter$count = 52842;
	#10 counter$count = 52843;
	#10 counter$count = 52844;
	#10 counter$count = 52845;
	#10 counter$count = 52846;
	#10 counter$count = 52847;
	#10 counter$count = 52848;
	#10 counter$count = 52849;
	#10 counter$count = 52850;
	#10 counter$count = 52851;
	#10 counter$count = 52852;
	#10 counter$count = 52853;
	#10 counter$count = 52854;
	#10 counter$count = 52855;
	#10 counter$count = 52856;
	#10 counter$count = 52857;
	#10 counter$count = 52858;
	#10 counter$count = 52859;
	#10 counter$count = 52860;
	#10 counter$count = 52861;
	#10 counter$count = 52862;
	#10 counter$count = 52863;
	#10 counter$count = 52864;
	#10 counter$count = 52865;
	#10 counter$count = 52866;
	#10 counter$count = 52867;
	#10 counter$count = 52868;
	#10 counter$count = 52869;
	#10 counter$count = 52870;
	#10 counter$count = 52871;
	#10 counter$count = 52872;
	#10 counter$count = 52873;
	#10 counter$count = 52874;
	#10 counter$count = 52875;
	#10 counter$count = 52876;
	#10 counter$count = 52877;
	#10 counter$count = 52878;
	#10 counter$count = 52879;
	#10 counter$count = 52880;
	#10 counter$count = 52881;
	#10 counter$count = 52882;
	#10 counter$count = 52883;
	#10 counter$count = 52884;
	#10 counter$count = 52885;
	#10 counter$count = 52886;
	#10 counter$count = 52887;
	#10 counter$count = 52888;
	#10 counter$count = 52889;
	#10 counter$count = 52890;
	#10 counter$count = 52891;
	#10 counter$count = 52892;
	#10 counter$count = 52893;
	#10 counter$count = 52894;
	#10 counter$count = 52895;
	#10 counter$count = 52896;
	#10 counter$count = 52897;
	#10 counter$count = 52898;
	#10 counter$count = 52899;
	#10 counter$count = 52900;
	#10 counter$count = 52901;
	#10 counter$count = 52902;
	#10 counter$count = 52903;
	#10 counter$count = 52904;
	#10 counter$count = 52905;
	#10 counter$count = 52906;
	#10 counter$count = 52907;
	#10 counter$count = 52908;
	#10 counter$count = 52909;
	#10 counter$count = 52910;
	#10 counter$count = 52911;
	#10 counter$count = 52912;
	#10 counter$count = 52913;
	#10 counter$count = 52914;
	#10 counter$count = 52915;
	#10 counter$count = 52916;
	#10 counter$count = 52917;
	#10 counter$count = 52918;
	#10 counter$count = 52919;
	#10 counter$count = 52920;
	#10 counter$count = 52921;
	#10 counter$count = 52922;
	#10 counter$count = 52923;
	#10 counter$count = 52924;
	#10 counter$count = 52925;
	#10 counter$count = 52926;
	#10 counter$count = 52927;
	#10 counter$count = 52928;
	#10 counter$count = 52929;
	#10 counter$count = 52930;
	#10 counter$count = 52931;
	#10 counter$count = 52932;
	#10 counter$count = 52933;
	#10 counter$count = 52934;
	#10 counter$count = 52935;
	#10 counter$count = 52936;
	#10 counter$count = 52937;
	#10 counter$count = 52938;
	#10 counter$count = 52939;
	#10 counter$count = 52940;
	#10 counter$count = 52941;
	#10 counter$count = 52942;
	#10 counter$count = 52943;
	#10 counter$count = 52944;
	#10 counter$count = 52945;
	#10 counter$count = 52946;
	#10 counter$count = 52947;
	#10 counter$count = 52948;
	#10 counter$count = 52949;
	#10 counter$count = 52950;
	#10 counter$count = 52951;
	#10 counter$count = 52952;
	#10 counter$count = 52953;
	#10 counter$count = 52954;
	#10 counter$count = 52955;
	#10 counter$count = 52956;
	#10 counter$count = 52957;
	#10 counter$count = 52958;
	#10 counter$count = 52959;
	#10 counter$count = 52960;
	#10 counter$count = 52961;
	#10 counter$count = 52962;
	#10 counter$count = 52963;
	#10 counter$count = 52964;
	#10 counter$count = 52965;
	#10 counter$count = 52966;
	#10 counter$count = 52967;
	#10 counter$count = 52968;
	#10 counter$count = 52969;
	#10 counter$count = 52970;
	#10 counter$count = 52971;
	#10 counter$count = 52972;
	#10 counter$count = 52973;
	#10 counter$count = 52974;
	#10 counter$count = 52975;
	#10 counter$count = 52976;
	#10 counter$count = 52977;
	#10 counter$count = 52978;
	#10 counter$count = 52979;
	#10 counter$count = 52980;
	#10 counter$count = 52981;
	#10 counter$count = 52982;
	#10 counter$count = 52983;
	#10 counter$count = 52984;
	#10 counter$count = 52985;
	#10 counter$count = 52986;
	#10 counter$count = 52987;
	#10 counter$count = 52988;
	#10 counter$count = 52989;
	#10 counter$count = 52990;
	#10 counter$count = 52991;
	#10 counter$count = 52992;
	#10 counter$count = 52993;
	#10 counter$count = 52994;
	#10 counter$count = 52995;
	#10 counter$count = 52996;
	#10 counter$count = 52997;
	#10 counter$count = 52998;
	#10 counter$count = 52999;
	#10 counter$count = 53000;
	#10 counter$count = 53001;
	#10 counter$count = 53002;
	#10 counter$count = 53003;
	#10 counter$count = 53004;
	#10 counter$count = 53005;
	#10 counter$count = 53006;
	#10 counter$count = 53007;
	#10 counter$count = 53008;
	#10 counter$count = 53009;
	#10 counter$count = 53010;
	#10 counter$count = 53011;
	#10 counter$count = 53012;
	#10 counter$count = 53013;
	#10 counter$count = 53014;
	#10 counter$count = 53015;
	#10 counter$count = 53016;
	#10 counter$count = 53017;
	#10 counter$count = 53018;
	#10 counter$count = 53019;
	#10 counter$count = 53020;
	#10 counter$count = 53021;
	#10 counter$count = 53022;
	#10 counter$count = 53023;
	#10 counter$count = 53024;
	#10 counter$count = 53025;
	#10 counter$count = 53026;
	#10 counter$count = 53027;
	#10 counter$count = 53028;
	#10 counter$count = 53029;
	#10 counter$count = 53030;
	#10 counter$count = 53031;
	#10 counter$count = 53032;
	#10 counter$count = 53033;
	#10 counter$count = 53034;
	#10 counter$count = 53035;
	#10 counter$count = 53036;
	#10 counter$count = 53037;
	#10 counter$count = 53038;
	#10 counter$count = 53039;
	#10 counter$count = 53040;
	#10 counter$count = 53041;
	#10 counter$count = 53042;
	#10 counter$count = 53043;
	#10 counter$count = 53044;
	#10 counter$count = 53045;
	#10 counter$count = 53046;
	#10 counter$count = 53047;
	#10 counter$count = 53048;
	#10 counter$count = 53049;
	#10 counter$count = 53050;
	#10 counter$count = 53051;
	#10 counter$count = 53052;
	#10 counter$count = 53053;
	#10 counter$count = 53054;
	#10 counter$count = 53055;
	#10 counter$count = 53056;
	#10 counter$count = 53057;
	#10 counter$count = 53058;
	#10 counter$count = 53059;
	#10 counter$count = 53060;
	#10 counter$count = 53061;
	#10 counter$count = 53062;
	#10 counter$count = 53063;
	#10 counter$count = 53064;
	#10 counter$count = 53065;
	#10 counter$count = 53066;
	#10 counter$count = 53067;
	#10 counter$count = 53068;
	#10 counter$count = 53069;
	#10 counter$count = 53070;
	#10 counter$count = 53071;
	#10 counter$count = 53072;
	#10 counter$count = 53073;
	#10 counter$count = 53074;
	#10 counter$count = 53075;
	#10 counter$count = 53076;
	#10 counter$count = 53077;
	#10 counter$count = 53078;
	#10 counter$count = 53079;
	#10 counter$count = 53080;
	#10 counter$count = 53081;
	#10 counter$count = 53082;
	#10 counter$count = 53083;
	#10 counter$count = 53084;
	#10 counter$count = 53085;
	#10 counter$count = 53086;
	#10 counter$count = 53087;
	#10 counter$count = 53088;
	#10 counter$count = 53089;
	#10 counter$count = 53090;
	#10 counter$count = 53091;
	#10 counter$count = 53092;
	#10 counter$count = 53093;
	#10 counter$count = 53094;
	#10 counter$count = 53095;
	#10 counter$count = 53096;
	#10 counter$count = 53097;
	#10 counter$count = 53098;
	#10 counter$count = 53099;
	#10 counter$count = 53100;
	#10 counter$count = 53101;
	#10 counter$count = 53102;
	#10 counter$count = 53103;
	#10 counter$count = 53104;
	#10 counter$count = 53105;
	#10 counter$count = 53106;
	#10 counter$count = 53107;
	#10 counter$count = 53108;
	#10 counter$count = 53109;
	#10 counter$count = 53110;
	#10 counter$count = 53111;
	#10 counter$count = 53112;
	#10 counter$count = 53113;
	#10 counter$count = 53114;
	#10 counter$count = 53115;
	#10 counter$count = 53116;
	#10 counter$count = 53117;
	#10 counter$count = 53118;
	#10 counter$count = 53119;
	#10 counter$count = 53120;
	#10 counter$count = 53121;
	#10 counter$count = 53122;
	#10 counter$count = 53123;
	#10 counter$count = 53124;
	#10 counter$count = 53125;
	#10 counter$count = 53126;
	#10 counter$count = 53127;
	#10 counter$count = 53128;
	#10 counter$count = 53129;
	#10 counter$count = 53130;
	#10 counter$count = 53131;
	#10 counter$count = 53132;
	#10 counter$count = 53133;
	#10 counter$count = 53134;
	#10 counter$count = 53135;
	#10 counter$count = 53136;
	#10 counter$count = 53137;
	#10 counter$count = 53138;
	#10 counter$count = 53139;
	#10 counter$count = 53140;
	#10 counter$count = 53141;
	#10 counter$count = 53142;
	#10 counter$count = 53143;
	#10 counter$count = 53144;
	#10 counter$count = 53145;
	#10 counter$count = 53146;
	#10 counter$count = 53147;
	#10 counter$count = 53148;
	#10 counter$count = 53149;
	#10 counter$count = 53150;
	#10 counter$count = 53151;
	#10 counter$count = 53152;
	#10 counter$count = 53153;
	#10 counter$count = 53154;
	#10 counter$count = 53155;
	#10 counter$count = 53156;
	#10 counter$count = 53157;
	#10 counter$count = 53158;
	#10 counter$count = 53159;
	#10 counter$count = 53160;
	#10 counter$count = 53161;
	#10 counter$count = 53162;
	#10 counter$count = 53163;
	#10 counter$count = 53164;
	#10 counter$count = 53165;
	#10 counter$count = 53166;
	#10 counter$count = 53167;
	#10 counter$count = 53168;
	#10 counter$count = 53169;
	#10 counter$count = 53170;
	#10 counter$count = 53171;
	#10 counter$count = 53172;
	#10 counter$count = 53173;
	#10 counter$count = 53174;
	#10 counter$count = 53175;
	#10 counter$count = 53176;
	#10 counter$count = 53177;
	#10 counter$count = 53178;
	#10 counter$count = 53179;
	#10 counter$count = 53180;
	#10 counter$count = 53181;
	#10 counter$count = 53182;
	#10 counter$count = 53183;
	#10 counter$count = 53184;
	#10 counter$count = 53185;
	#10 counter$count = 53186;
	#10 counter$count = 53187;
	#10 counter$count = 53188;
	#10 counter$count = 53189;
	#10 counter$count = 53190;
	#10 counter$count = 53191;
	#10 counter$count = 53192;
	#10 counter$count = 53193;
	#10 counter$count = 53194;
	#10 counter$count = 53195;
	#10 counter$count = 53196;
	#10 counter$count = 53197;
	#10 counter$count = 53198;
	#10 counter$count = 53199;
	#10 counter$count = 53200;
	#10 counter$count = 53201;
	#10 counter$count = 53202;
	#10 counter$count = 53203;
	#10 counter$count = 53204;
	#10 counter$count = 53205;
	#10 counter$count = 53206;
	#10 counter$count = 53207;
	#10 counter$count = 53208;
	#10 counter$count = 53209;
	#10 counter$count = 53210;
	#10 counter$count = 53211;
	#10 counter$count = 53212;
	#10 counter$count = 53213;
	#10 counter$count = 53214;
	#10 counter$count = 53215;
	#10 counter$count = 53216;
	#10 counter$count = 53217;
	#10 counter$count = 53218;
	#10 counter$count = 53219;
	#10 counter$count = 53220;
	#10 counter$count = 53221;
	#10 counter$count = 53222;
	#10 counter$count = 53223;
	#10 counter$count = 53224;
	#10 counter$count = 53225;
	#10 counter$count = 53226;
	#10 counter$count = 53227;
	#10 counter$count = 53228;
	#10 counter$count = 53229;
	#10 counter$count = 53230;
	#10 counter$count = 53231;
	#10 counter$count = 53232;
	#10 counter$count = 53233;
	#10 counter$count = 53234;
	#10 counter$count = 53235;
	#10 counter$count = 53236;
	#10 counter$count = 53237;
	#10 counter$count = 53238;
	#10 counter$count = 53239;
	#10 counter$count = 53240;
	#10 counter$count = 53241;
	#10 counter$count = 53242;
	#10 counter$count = 53243;
	#10 counter$count = 53244;
	#10 counter$count = 53245;
	#10 counter$count = 53246;
	#10 counter$count = 53247;
	#10 counter$count = 53248;
	#10 counter$count = 53249;
	#10 counter$count = 53250;
	#10 counter$count = 53251;
	#10 counter$count = 53252;
	#10 counter$count = 53253;
	#10 counter$count = 53254;
	#10 counter$count = 53255;
	#10 counter$count = 53256;
	#10 counter$count = 53257;
	#10 counter$count = 53258;
	#10 counter$count = 53259;
	#10 counter$count = 53260;
	#10 counter$count = 53261;
	#10 counter$count = 53262;
	#10 counter$count = 53263;
	#10 counter$count = 53264;
	#10 counter$count = 53265;
	#10 counter$count = 53266;
	#10 counter$count = 53267;
	#10 counter$count = 53268;
	#10 counter$count = 53269;
	#10 counter$count = 53270;
	#10 counter$count = 53271;
	#10 counter$count = 53272;
	#10 counter$count = 53273;
	#10 counter$count = 53274;
	#10 counter$count = 53275;
	#10 counter$count = 53276;
	#10 counter$count = 53277;
	#10 counter$count = 53278;
	#10 counter$count = 53279;
	#10 counter$count = 53280;
	#10 counter$count = 53281;
	#10 counter$count = 53282;
	#10 counter$count = 53283;
	#10 counter$count = 53284;
	#10 counter$count = 53285;
	#10 counter$count = 53286;
	#10 counter$count = 53287;
	#10 counter$count = 53288;
	#10 counter$count = 53289;
	#10 counter$count = 53290;
	#10 counter$count = 53291;
	#10 counter$count = 53292;
	#10 counter$count = 53293;
	#10 counter$count = 53294;
	#10 counter$count = 53295;
	#10 counter$count = 53296;
	#10 counter$count = 53297;
	#10 counter$count = 53298;
	#10 counter$count = 53299;
	#10 counter$count = 53300;
	#10 counter$count = 53301;
	#10 counter$count = 53302;
	#10 counter$count = 53303;
	#10 counter$count = 53304;
	#10 counter$count = 53305;
	#10 counter$count = 53306;
	#10 counter$count = 53307;
	#10 counter$count = 53308;
	#10 counter$count = 53309;
	#10 counter$count = 53310;
	#10 counter$count = 53311;
	#10 counter$count = 53312;
	#10 counter$count = 53313;
	#10 counter$count = 53314;
	#10 counter$count = 53315;
	#10 counter$count = 53316;
	#10 counter$count = 53317;
	#10 counter$count = 53318;
	#10 counter$count = 53319;
	#10 counter$count = 53320;
	#10 counter$count = 53321;
	#10 counter$count = 53322;
	#10 counter$count = 53323;
	#10 counter$count = 53324;
	#10 counter$count = 53325;
	#10 counter$count = 53326;
	#10 counter$count = 53327;
	#10 counter$count = 53328;
	#10 counter$count = 53329;
	#10 counter$count = 53330;
	#10 counter$count = 53331;
	#10 counter$count = 53332;
	#10 counter$count = 53333;
	#10 counter$count = 53334;
	#10 counter$count = 53335;
	#10 counter$count = 53336;
	#10 counter$count = 53337;
	#10 counter$count = 53338;
	#10 counter$count = 53339;
	#10 counter$count = 53340;
	#10 counter$count = 53341;
	#10 counter$count = 53342;
	#10 counter$count = 53343;
	#10 counter$count = 53344;
	#10 counter$count = 53345;
	#10 counter$count = 53346;
	#10 counter$count = 53347;
	#10 counter$count = 53348;
	#10 counter$count = 53349;
	#10 counter$count = 53350;
	#10 counter$count = 53351;
	#10 counter$count = 53352;
	#10 counter$count = 53353;
	#10 counter$count = 53354;
	#10 counter$count = 53355;
	#10 counter$count = 53356;
	#10 counter$count = 53357;
	#10 counter$count = 53358;
	#10 counter$count = 53359;
	#10 counter$count = 53360;
	#10 counter$count = 53361;
	#10 counter$count = 53362;
	#10 counter$count = 53363;
	#10 counter$count = 53364;
	#10 counter$count = 53365;
	#10 counter$count = 53366;
	#10 counter$count = 53367;
	#10 counter$count = 53368;
	#10 counter$count = 53369;
	#10 counter$count = 53370;
	#10 counter$count = 53371;
	#10 counter$count = 53372;
	#10 counter$count = 53373;
	#10 counter$count = 53374;
	#10 counter$count = 53375;
	#10 counter$count = 53376;
	#10 counter$count = 53377;
	#10 counter$count = 53378;
	#10 counter$count = 53379;
	#10 counter$count = 53380;
	#10 counter$count = 53381;
	#10 counter$count = 53382;
	#10 counter$count = 53383;
	#10 counter$count = 53384;
	#10 counter$count = 53385;
	#10 counter$count = 53386;
	#10 counter$count = 53387;
	#10 counter$count = 53388;
	#10 counter$count = 53389;
	#10 counter$count = 53390;
	#10 counter$count = 53391;
	#10 counter$count = 53392;
	#10 counter$count = 53393;
	#10 counter$count = 53394;
	#10 counter$count = 53395;
	#10 counter$count = 53396;
	#10 counter$count = 53397;
	#10 counter$count = 53398;
	#10 counter$count = 53399;
	#10 counter$count = 53400;
	#10 counter$count = 53401;
	#10 counter$count = 53402;
	#10 counter$count = 53403;
	#10 counter$count = 53404;
	#10 counter$count = 53405;
	#10 counter$count = 53406;
	#10 counter$count = 53407;
	#10 counter$count = 53408;
	#10 counter$count = 53409;
	#10 counter$count = 53410;
	#10 counter$count = 53411;
	#10 counter$count = 53412;
	#10 counter$count = 53413;
	#10 counter$count = 53414;
	#10 counter$count = 53415;
	#10 counter$count = 53416;
	#10 counter$count = 53417;
	#10 counter$count = 53418;
	#10 counter$count = 53419;
	#10 counter$count = 53420;
	#10 counter$count = 53421;
	#10 counter$count = 53422;
	#10 counter$count = 53423;
	#10 counter$count = 53424;
	#10 counter$count = 53425;
	#10 counter$count = 53426;
	#10 counter$count = 53427;
	#10 counter$count = 53428;
	#10 counter$count = 53429;
	#10 counter$count = 53430;
	#10 counter$count = 53431;
	#10 counter$count = 53432;
	#10 counter$count = 53433;
	#10 counter$count = 53434;
	#10 counter$count = 53435;
	#10 counter$count = 53436;
	#10 counter$count = 53437;
	#10 counter$count = 53438;
	#10 counter$count = 53439;
	#10 counter$count = 53440;
	#10 counter$count = 53441;
	#10 counter$count = 53442;
	#10 counter$count = 53443;
	#10 counter$count = 53444;
	#10 counter$count = 53445;
	#10 counter$count = 53446;
	#10 counter$count = 53447;
	#10 counter$count = 53448;
	#10 counter$count = 53449;
	#10 counter$count = 53450;
	#10 counter$count = 53451;
	#10 counter$count = 53452;
	#10 counter$count = 53453;
	#10 counter$count = 53454;
	#10 counter$count = 53455;
	#10 counter$count = 53456;
	#10 counter$count = 53457;
	#10 counter$count = 53458;
	#10 counter$count = 53459;
	#10 counter$count = 53460;
	#10 counter$count = 53461;
	#10 counter$count = 53462;
	#10 counter$count = 53463;
	#10 counter$count = 53464;
	#10 counter$count = 53465;
	#10 counter$count = 53466;
	#10 counter$count = 53467;
	#10 counter$count = 53468;
	#10 counter$count = 53469;
	#10 counter$count = 53470;
	#10 counter$count = 53471;
	#10 counter$count = 53472;
	#10 counter$count = 53473;
	#10 counter$count = 53474;
	#10 counter$count = 53475;
	#10 counter$count = 53476;
	#10 counter$count = 53477;
	#10 counter$count = 53478;
	#10 counter$count = 53479;
	#10 counter$count = 53480;
	#10 counter$count = 53481;
	#10 counter$count = 53482;
	#10 counter$count = 53483;
	#10 counter$count = 53484;
	#10 counter$count = 53485;
	#10 counter$count = 53486;
	#10 counter$count = 53487;
	#10 counter$count = 53488;
	#10 counter$count = 53489;
	#10 counter$count = 53490;
	#10 counter$count = 53491;
	#10 counter$count = 53492;
	#10 counter$count = 53493;
	#10 counter$count = 53494;
	#10 counter$count = 53495;
	#10 counter$count = 53496;
	#10 counter$count = 53497;
	#10 counter$count = 53498;
	#10 counter$count = 53499;
	#10 counter$count = 53500;
	#10 counter$count = 53501;
	#10 counter$count = 53502;
	#10 counter$count = 53503;
	#10 counter$count = 53504;
	#10 counter$count = 53505;
	#10 counter$count = 53506;
	#10 counter$count = 53507;
	#10 counter$count = 53508;
	#10 counter$count = 53509;
	#10 counter$count = 53510;
	#10 counter$count = 53511;
	#10 counter$count = 53512;
	#10 counter$count = 53513;
	#10 counter$count = 53514;
	#10 counter$count = 53515;
	#10 counter$count = 53516;
	#10 counter$count = 53517;
	#10 counter$count = 53518;
	#10 counter$count = 53519;
	#10 counter$count = 53520;
	#10 counter$count = 53521;
	#10 counter$count = 53522;
	#10 counter$count = 53523;
	#10 counter$count = 53524;
	#10 counter$count = 53525;
	#10 counter$count = 53526;
	#10 counter$count = 53527;
	#10 counter$count = 53528;
	#10 counter$count = 53529;
	#10 counter$count = 53530;
	#10 counter$count = 53531;
	#10 counter$count = 53532;
	#10 counter$count = 53533;
	#10 counter$count = 53534;
	#10 counter$count = 53535;
	#10 counter$count = 53536;
	#10 counter$count = 53537;
	#10 counter$count = 53538;
	#10 counter$count = 53539;
	#10 counter$count = 53540;
	#10 counter$count = 53541;
	#10 counter$count = 53542;
	#10 counter$count = 53543;
	#10 counter$count = 53544;
	#10 counter$count = 53545;
	#10 counter$count = 53546;
	#10 counter$count = 53547;
	#10 counter$count = 53548;
	#10 counter$count = 53549;
	#10 counter$count = 53550;
	#10 counter$count = 53551;
	#10 counter$count = 53552;
	#10 counter$count = 53553;
	#10 counter$count = 53554;
	#10 counter$count = 53555;
	#10 counter$count = 53556;
	#10 counter$count = 53557;
	#10 counter$count = 53558;
	#10 counter$count = 53559;
	#10 counter$count = 53560;
	#10 counter$count = 53561;
	#10 counter$count = 53562;
	#10 counter$count = 53563;
	#10 counter$count = 53564;
	#10 counter$count = 53565;
	#10 counter$count = 53566;
	#10 counter$count = 53567;
	#10 counter$count = 53568;
	#10 counter$count = 53569;
	#10 counter$count = 53570;
	#10 counter$count = 53571;
	#10 counter$count = 53572;
	#10 counter$count = 53573;
	#10 counter$count = 53574;
	#10 counter$count = 53575;
	#10 counter$count = 53576;
	#10 counter$count = 53577;
	#10 counter$count = 53578;
	#10 counter$count = 53579;
	#10 counter$count = 53580;
	#10 counter$count = 53581;
	#10 counter$count = 53582;
	#10 counter$count = 53583;
	#10 counter$count = 53584;
	#10 counter$count = 53585;
	#10 counter$count = 53586;
	#10 counter$count = 53587;
	#10 counter$count = 53588;
	#10 counter$count = 53589;
	#10 counter$count = 53590;
	#10 counter$count = 53591;
	#10 counter$count = 53592;
	#10 counter$count = 53593;
	#10 counter$count = 53594;
	#10 counter$count = 53595;
	#10 counter$count = 53596;
	#10 counter$count = 53597;
	#10 counter$count = 53598;
	#10 counter$count = 53599;
	#10 counter$count = 53600;
	#10 counter$count = 53601;
	#10 counter$count = 53602;
	#10 counter$count = 53603;
	#10 counter$count = 53604;
	#10 counter$count = 53605;
	#10 counter$count = 53606;
	#10 counter$count = 53607;
	#10 counter$count = 53608;
	#10 counter$count = 53609;
	#10 counter$count = 53610;
	#10 counter$count = 53611;
	#10 counter$count = 53612;
	#10 counter$count = 53613;
	#10 counter$count = 53614;
	#10 counter$count = 53615;
	#10 counter$count = 53616;
	#10 counter$count = 53617;
	#10 counter$count = 53618;
	#10 counter$count = 53619;
	#10 counter$count = 53620;
	#10 counter$count = 53621;
	#10 counter$count = 53622;
	#10 counter$count = 53623;
	#10 counter$count = 53624;
	#10 counter$count = 53625;
	#10 counter$count = 53626;
	#10 counter$count = 53627;
	#10 counter$count = 53628;
	#10 counter$count = 53629;
	#10 counter$count = 53630;
	#10 counter$count = 53631;
	#10 counter$count = 53632;
	#10 counter$count = 53633;
	#10 counter$count = 53634;
	#10 counter$count = 53635;
	#10 counter$count = 53636;
	#10 counter$count = 53637;
	#10 counter$count = 53638;
	#10 counter$count = 53639;
	#10 counter$count = 53640;
	#10 counter$count = 53641;
	#10 counter$count = 53642;
	#10 counter$count = 53643;
	#10 counter$count = 53644;
	#10 counter$count = 53645;
	#10 counter$count = 53646;
	#10 counter$count = 53647;
	#10 counter$count = 53648;
	#10 counter$count = 53649;
	#10 counter$count = 53650;
	#10 counter$count = 53651;
	#10 counter$count = 53652;
	#10 counter$count = 53653;
	#10 counter$count = 53654;
	#10 counter$count = 53655;
	#10 counter$count = 53656;
	#10 counter$count = 53657;
	#10 counter$count = 53658;
	#10 counter$count = 53659;
	#10 counter$count = 53660;
	#10 counter$count = 53661;
	#10 counter$count = 53662;
	#10 counter$count = 53663;
	#10 counter$count = 53664;
	#10 counter$count = 53665;
	#10 counter$count = 53666;
	#10 counter$count = 53667;
	#10 counter$count = 53668;
	#10 counter$count = 53669;
	#10 counter$count = 53670;
	#10 counter$count = 53671;
	#10 counter$count = 53672;
	#10 counter$count = 53673;
	#10 counter$count = 53674;
	#10 counter$count = 53675;
	#10 counter$count = 53676;
	#10 counter$count = 53677;
	#10 counter$count = 53678;
	#10 counter$count = 53679;
	#10 counter$count = 53680;
	#10 counter$count = 53681;
	#10 counter$count = 53682;
	#10 counter$count = 53683;
	#10 counter$count = 53684;
	#10 counter$count = 53685;
	#10 counter$count = 53686;
	#10 counter$count = 53687;
	#10 counter$count = 53688;
	#10 counter$count = 53689;
	#10 counter$count = 53690;
	#10 counter$count = 53691;
	#10 counter$count = 53692;
	#10 counter$count = 53693;
	#10 counter$count = 53694;
	#10 counter$count = 53695;
	#10 counter$count = 53696;
	#10 counter$count = 53697;
	#10 counter$count = 53698;
	#10 counter$count = 53699;
	#10 counter$count = 53700;
	#10 counter$count = 53701;
	#10 counter$count = 53702;
	#10 counter$count = 53703;
	#10 counter$count = 53704;
	#10 counter$count = 53705;
	#10 counter$count = 53706;
	#10 counter$count = 53707;
	#10 counter$count = 53708;
	#10 counter$count = 53709;
	#10 counter$count = 53710;
	#10 counter$count = 53711;
	#10 counter$count = 53712;
	#10 counter$count = 53713;
	#10 counter$count = 53714;
	#10 counter$count = 53715;
	#10 counter$count = 53716;
	#10 counter$count = 53717;
	#10 counter$count = 53718;
	#10 counter$count = 53719;
	#10 counter$count = 53720;
	#10 counter$count = 53721;
	#10 counter$count = 53722;
	#10 counter$count = 53723;
	#10 counter$count = 53724;
	#10 counter$count = 53725;
	#10 counter$count = 53726;
	#10 counter$count = 53727;
	#10 counter$count = 53728;
	#10 counter$count = 53729;
	#10 counter$count = 53730;
	#10 counter$count = 53731;
	#10 counter$count = 53732;
	#10 counter$count = 53733;
	#10 counter$count = 53734;
	#10 counter$count = 53735;
	#10 counter$count = 53736;
	#10 counter$count = 53737;
	#10 counter$count = 53738;
	#10 counter$count = 53739;
	#10 counter$count = 53740;
	#10 counter$count = 53741;
	#10 counter$count = 53742;
	#10 counter$count = 53743;
	#10 counter$count = 53744;
	#10 counter$count = 53745;
	#10 counter$count = 53746;
	#10 counter$count = 53747;
	#10 counter$count = 53748;
	#10 counter$count = 53749;
	#10 counter$count = 53750;
	#10 counter$count = 53751;
	#10 counter$count = 53752;
	#10 counter$count = 53753;
	#10 counter$count = 53754;
	#10 counter$count = 53755;
	#10 counter$count = 53756;
	#10 counter$count = 53757;
	#10 counter$count = 53758;
	#10 counter$count = 53759;
	#10 counter$count = 53760;
	#10 counter$count = 53761;
	#10 counter$count = 53762;
	#10 counter$count = 53763;
	#10 counter$count = 53764;
	#10 counter$count = 53765;
	#10 counter$count = 53766;
	#10 counter$count = 53767;
	#10 counter$count = 53768;
	#10 counter$count = 53769;
	#10 counter$count = 53770;
	#10 counter$count = 53771;
	#10 counter$count = 53772;
	#10 counter$count = 53773;
	#10 counter$count = 53774;
	#10 counter$count = 53775;
	#10 counter$count = 53776;
	#10 counter$count = 53777;
	#10 counter$count = 53778;
	#10 counter$count = 53779;
	#10 counter$count = 53780;
	#10 counter$count = 53781;
	#10 counter$count = 53782;
	#10 counter$count = 53783;
	#10 counter$count = 53784;
	#10 counter$count = 53785;
	#10 counter$count = 53786;
	#10 counter$count = 53787;
	#10 counter$count = 53788;
	#10 counter$count = 53789;
	#10 counter$count = 53790;
	#10 counter$count = 53791;
	#10 counter$count = 53792;
	#10 counter$count = 53793;
	#10 counter$count = 53794;
	#10 counter$count = 53795;
	#10 counter$count = 53796;
	#10 counter$count = 53797;
	#10 counter$count = 53798;
	#10 counter$count = 53799;
	#10 counter$count = 53800;
	#10 counter$count = 53801;
	#10 counter$count = 53802;
	#10 counter$count = 53803;
	#10 counter$count = 53804;
	#10 counter$count = 53805;
	#10 counter$count = 53806;
	#10 counter$count = 53807;
	#10 counter$count = 53808;
	#10 counter$count = 53809;
	#10 counter$count = 53810;
	#10 counter$count = 53811;
	#10 counter$count = 53812;
	#10 counter$count = 53813;
	#10 counter$count = 53814;
	#10 counter$count = 53815;
	#10 counter$count = 53816;
	#10 counter$count = 53817;
	#10 counter$count = 53818;
	#10 counter$count = 53819;
	#10 counter$count = 53820;
	#10 counter$count = 53821;
	#10 counter$count = 53822;
	#10 counter$count = 53823;
	#10 counter$count = 53824;
	#10 counter$count = 53825;
	#10 counter$count = 53826;
	#10 counter$count = 53827;
	#10 counter$count = 53828;
	#10 counter$count = 53829;
	#10 counter$count = 53830;
	#10 counter$count = 53831;
	#10 counter$count = 53832;
	#10 counter$count = 53833;
	#10 counter$count = 53834;
	#10 counter$count = 53835;
	#10 counter$count = 53836;
	#10 counter$count = 53837;
	#10 counter$count = 53838;
	#10 counter$count = 53839;
	#10 counter$count = 53840;
	#10 counter$count = 53841;
	#10 counter$count = 53842;
	#10 counter$count = 53843;
	#10 counter$count = 53844;
	#10 counter$count = 53845;
	#10 counter$count = 53846;
	#10 counter$count = 53847;
	#10 counter$count = 53848;
	#10 counter$count = 53849;
	#10 counter$count = 53850;
	#10 counter$count = 53851;
	#10 counter$count = 53852;
	#10 counter$count = 53853;
	#10 counter$count = 53854;
	#10 counter$count = 53855;
	#10 counter$count = 53856;
	#10 counter$count = 53857;
	#10 counter$count = 53858;
	#10 counter$count = 53859;
	#10 counter$count = 53860;
	#10 counter$count = 53861;
	#10 counter$count = 53862;
	#10 counter$count = 53863;
	#10 counter$count = 53864;
	#10 counter$count = 53865;
	#10 counter$count = 53866;
	#10 counter$count = 53867;
	#10 counter$count = 53868;
	#10 counter$count = 53869;
	#10 counter$count = 53870;
	#10 counter$count = 53871;
	#10 counter$count = 53872;
	#10 counter$count = 53873;
	#10 counter$count = 53874;
	#10 counter$count = 53875;
	#10 counter$count = 53876;
	#10 counter$count = 53877;
	#10 counter$count = 53878;
	#10 counter$count = 53879;
	#10 counter$count = 53880;
	#10 counter$count = 53881;
	#10 counter$count = 53882;
	#10 counter$count = 53883;
	#10 counter$count = 53884;
	#10 counter$count = 53885;
	#10 counter$count = 53886;
	#10 counter$count = 53887;
	#10 counter$count = 53888;
	#10 counter$count = 53889;
	#10 counter$count = 53890;
	#10 counter$count = 53891;
	#10 counter$count = 53892;
	#10 counter$count = 53893;
	#10 counter$count = 53894;
	#10 counter$count = 53895;
	#10 counter$count = 53896;
	#10 counter$count = 53897;
	#10 counter$count = 53898;
	#10 counter$count = 53899;
	#10 counter$count = 53900;
	#10 counter$count = 53901;
	#10 counter$count = 53902;
	#10 counter$count = 53903;
	#10 counter$count = 53904;
	#10 counter$count = 53905;
	#10 counter$count = 53906;
	#10 counter$count = 53907;
	#10 counter$count = 53908;
	#10 counter$count = 53909;
	#10 counter$count = 53910;
	#10 counter$count = 53911;
	#10 counter$count = 53912;
	#10 counter$count = 53913;
	#10 counter$count = 53914;
	#10 counter$count = 53915;
	#10 counter$count = 53916;
	#10 counter$count = 53917;
	#10 counter$count = 53918;
	#10 counter$count = 53919;
	#10 counter$count = 53920;
	#10 counter$count = 53921;
	#10 counter$count = 53922;
	#10 counter$count = 53923;
	#10 counter$count = 53924;
	#10 counter$count = 53925;
	#10 counter$count = 53926;
	#10 counter$count = 53927;
	#10 counter$count = 53928;
	#10 counter$count = 53929;
	#10 counter$count = 53930;
	#10 counter$count = 53931;
	#10 counter$count = 53932;
	#10 counter$count = 53933;
	#10 counter$count = 53934;
	#10 counter$count = 53935;
	#10 counter$count = 53936;
	#10 counter$count = 53937;
	#10 counter$count = 53938;
	#10 counter$count = 53939;
	#10 counter$count = 53940;
	#10 counter$count = 53941;
	#10 counter$count = 53942;
	#10 counter$count = 53943;
	#10 counter$count = 53944;
	#10 counter$count = 53945;
	#10 counter$count = 53946;
	#10 counter$count = 53947;
	#10 counter$count = 53948;
	#10 counter$count = 53949;
	#10 counter$count = 53950;
	#10 counter$count = 53951;
	#10 counter$count = 53952;
	#10 counter$count = 53953;
	#10 counter$count = 53954;
	#10 counter$count = 53955;
	#10 counter$count = 53956;
	#10 counter$count = 53957;
	#10 counter$count = 53958;
	#10 counter$count = 53959;
	#10 counter$count = 53960;
	#10 counter$count = 53961;
	#10 counter$count = 53962;
	#10 counter$count = 53963;
	#10 counter$count = 53964;
	#10 counter$count = 53965;
	#10 counter$count = 53966;
	#10 counter$count = 53967;
	#10 counter$count = 53968;
	#10 counter$count = 53969;
	#10 counter$count = 53970;
	#10 counter$count = 53971;
	#10 counter$count = 53972;
	#10 counter$count = 53973;
	#10 counter$count = 53974;
	#10 counter$count = 53975;
	#10 counter$count = 53976;
	#10 counter$count = 53977;
	#10 counter$count = 53978;
	#10 counter$count = 53979;
	#10 counter$count = 53980;
	#10 counter$count = 53981;
	#10 counter$count = 53982;
	#10 counter$count = 53983;
	#10 counter$count = 53984;
	#10 counter$count = 53985;
	#10 counter$count = 53986;
	#10 counter$count = 53987;
	#10 counter$count = 53988;
	#10 counter$count = 53989;
	#10 counter$count = 53990;
	#10 counter$count = 53991;
	#10 counter$count = 53992;
	#10 counter$count = 53993;
	#10 counter$count = 53994;
	#10 counter$count = 53995;
	#10 counter$count = 53996;
	#10 counter$count = 53997;
	#10 counter$count = 53998;
	#10 counter$count = 53999;
	#10 counter$count = 54000;
	#10 counter$count = 54001;
	#10 counter$count = 54002;
	#10 counter$count = 54003;
	#10 counter$count = 54004;
	#10 counter$count = 54005;
	#10 counter$count = 54006;
	#10 counter$count = 54007;
	#10 counter$count = 54008;
	#10 counter$count = 54009;
	#10 counter$count = 54010;
	#10 counter$count = 54011;
	#10 counter$count = 54012;
	#10 counter$count = 54013;
	#10 counter$count = 54014;
	#10 counter$count = 54015;
	#10 counter$count = 54016;
	#10 counter$count = 54017;
	#10 counter$count = 54018;
	#10 counter$count = 54019;
	#10 counter$count = 54020;
	#10 counter$count = 54021;
	#10 counter$count = 54022;
	#10 counter$count = 54023;
	#10 counter$count = 54024;
	#10 counter$count = 54025;
	#10 counter$count = 54026;
	#10 counter$count = 54027;
	#10 counter$count = 54028;
	#10 counter$count = 54029;
	#10 counter$count = 54030;
	#10 counter$count = 54031;
	#10 counter$count = 54032;
	#10 counter$count = 54033;
	#10 counter$count = 54034;
	#10 counter$count = 54035;
	#10 counter$count = 54036;
	#10 counter$count = 54037;
	#10 counter$count = 54038;
	#10 counter$count = 54039;
	#10 counter$count = 54040;
	#10 counter$count = 54041;
	#10 counter$count = 54042;
	#10 counter$count = 54043;
	#10 counter$count = 54044;
	#10 counter$count = 54045;
	#10 counter$count = 54046;
	#10 counter$count = 54047;
	#10 counter$count = 54048;
	#10 counter$count = 54049;
	#10 counter$count = 54050;
	#10 counter$count = 54051;
	#10 counter$count = 54052;
	#10 counter$count = 54053;
	#10 counter$count = 54054;
	#10 counter$count = 54055;
	#10 counter$count = 54056;
	#10 counter$count = 54057;
	#10 counter$count = 54058;
	#10 counter$count = 54059;
	#10 counter$count = 54060;
	#10 counter$count = 54061;
	#10 counter$count = 54062;
	#10 counter$count = 54063;
	#10 counter$count = 54064;
	#10 counter$count = 54065;
	#10 counter$count = 54066;
	#10 counter$count = 54067;
	#10 counter$count = 54068;
	#10 counter$count = 54069;
	#10 counter$count = 54070;
	#10 counter$count = 54071;
	#10 counter$count = 54072;
	#10 counter$count = 54073;
	#10 counter$count = 54074;
	#10 counter$count = 54075;
	#10 counter$count = 54076;
	#10 counter$count = 54077;
	#10 counter$count = 54078;
	#10 counter$count = 54079;
	#10 counter$count = 54080;
	#10 counter$count = 54081;
	#10 counter$count = 54082;
	#10 counter$count = 54083;
	#10 counter$count = 54084;
	#10 counter$count = 54085;
	#10 counter$count = 54086;
	#10 counter$count = 54087;
	#10 counter$count = 54088;
	#10 counter$count = 54089;
	#10 counter$count = 54090;
	#10 counter$count = 54091;
	#10 counter$count = 54092;
	#10 counter$count = 54093;
	#10 counter$count = 54094;
	#10 counter$count = 54095;
	#10 counter$count = 54096;
	#10 counter$count = 54097;
	#10 counter$count = 54098;
	#10 counter$count = 54099;
	#10 counter$count = 54100;
	#10 counter$count = 54101;
	#10 counter$count = 54102;
	#10 counter$count = 54103;
	#10 counter$count = 54104;
	#10 counter$count = 54105;
	#10 counter$count = 54106;
	#10 counter$count = 54107;
	#10 counter$count = 54108;
	#10 counter$count = 54109;
	#10 counter$count = 54110;
	#10 counter$count = 54111;
	#10 counter$count = 54112;
	#10 counter$count = 54113;
	#10 counter$count = 54114;
	#10 counter$count = 54115;
	#10 counter$count = 54116;
	#10 counter$count = 54117;
	#10 counter$count = 54118;
	#10 counter$count = 54119;
	#10 counter$count = 54120;
	#10 counter$count = 54121;
	#10 counter$count = 54122;
	#10 counter$count = 54123;
	#10 counter$count = 54124;
	#10 counter$count = 54125;
	#10 counter$count = 54126;
	#10 counter$count = 54127;
	#10 counter$count = 54128;
	#10 counter$count = 54129;
	#10 counter$count = 54130;
	#10 counter$count = 54131;
	#10 counter$count = 54132;
	#10 counter$count = 54133;
	#10 counter$count = 54134;
	#10 counter$count = 54135;
	#10 counter$count = 54136;
	#10 counter$count = 54137;
	#10 counter$count = 54138;
	#10 counter$count = 54139;
	#10 counter$count = 54140;
	#10 counter$count = 54141;
	#10 counter$count = 54142;
	#10 counter$count = 54143;
	#10 counter$count = 54144;
	#10 counter$count = 54145;
	#10 counter$count = 54146;
	#10 counter$count = 54147;
	#10 counter$count = 54148;
	#10 counter$count = 54149;
	#10 counter$count = 54150;
	#10 counter$count = 54151;
	#10 counter$count = 54152;
	#10 counter$count = 54153;
	#10 counter$count = 54154;
	#10 counter$count = 54155;
	#10 counter$count = 54156;
	#10 counter$count = 54157;
	#10 counter$count = 54158;
	#10 counter$count = 54159;
	#10 counter$count = 54160;
	#10 counter$count = 54161;
	#10 counter$count = 54162;
	#10 counter$count = 54163;
	#10 counter$count = 54164;
	#10 counter$count = 54165;
	#10 counter$count = 54166;
	#10 counter$count = 54167;
	#10 counter$count = 54168;
	#10 counter$count = 54169;
	#10 counter$count = 54170;
	#10 counter$count = 54171;
	#10 counter$count = 54172;
	#10 counter$count = 54173;
	#10 counter$count = 54174;
	#10 counter$count = 54175;
	#10 counter$count = 54176;
	#10 counter$count = 54177;
	#10 counter$count = 54178;
	#10 counter$count = 54179;
	#10 counter$count = 54180;
	#10 counter$count = 54181;
	#10 counter$count = 54182;
	#10 counter$count = 54183;
	#10 counter$count = 54184;
	#10 counter$count = 54185;
	#10 counter$count = 54186;
	#10 counter$count = 54187;
	#10 counter$count = 54188;
	#10 counter$count = 54189;
	#10 counter$count = 54190;
	#10 counter$count = 54191;
	#10 counter$count = 54192;
	#10 counter$count = 54193;
	#10 counter$count = 54194;
	#10 counter$count = 54195;
	#10 counter$count = 54196;
	#10 counter$count = 54197;
	#10 counter$count = 54198;
	#10 counter$count = 54199;
	#10 counter$count = 54200;
	#10 counter$count = 54201;
	#10 counter$count = 54202;
	#10 counter$count = 54203;
	#10 counter$count = 54204;
	#10 counter$count = 54205;
	#10 counter$count = 54206;
	#10 counter$count = 54207;
	#10 counter$count = 54208;
	#10 counter$count = 54209;
	#10 counter$count = 54210;
	#10 counter$count = 54211;
	#10 counter$count = 54212;
	#10 counter$count = 54213;
	#10 counter$count = 54214;
	#10 counter$count = 54215;
	#10 counter$count = 54216;
	#10 counter$count = 54217;
	#10 counter$count = 54218;
	#10 counter$count = 54219;
	#10 counter$count = 54220;
	#10 counter$count = 54221;
	#10 counter$count = 54222;
	#10 counter$count = 54223;
	#10 counter$count = 54224;
	#10 counter$count = 54225;
	#10 counter$count = 54226;
	#10 counter$count = 54227;
	#10 counter$count = 54228;
	#10 counter$count = 54229;
	#10 counter$count = 54230;
	#10 counter$count = 54231;
	#10 counter$count = 54232;
	#10 counter$count = 54233;
	#10 counter$count = 54234;
	#10 counter$count = 54235;
	#10 counter$count = 54236;
	#10 counter$count = 54237;
	#10 counter$count = 54238;
	#10 counter$count = 54239;
	#10 counter$count = 54240;
	#10 counter$count = 54241;
	#10 counter$count = 54242;
	#10 counter$count = 54243;
	#10 counter$count = 54244;
	#10 counter$count = 54245;
	#10 counter$count = 54246;
	#10 counter$count = 54247;
	#10 counter$count = 54248;
	#10 counter$count = 54249;
	#10 counter$count = 54250;
	#10 counter$count = 54251;
	#10 counter$count = 54252;
	#10 counter$count = 54253;
	#10 counter$count = 54254;
	#10 counter$count = 54255;
	#10 counter$count = 54256;
	#10 counter$count = 54257;
	#10 counter$count = 54258;
	#10 counter$count = 54259;
	#10 counter$count = 54260;
	#10 counter$count = 54261;
	#10 counter$count = 54262;
	#10 counter$count = 54263;
	#10 counter$count = 54264;
	#10 counter$count = 54265;
	#10 counter$count = 54266;
	#10 counter$count = 54267;
	#10 counter$count = 54268;
	#10 counter$count = 54269;
	#10 counter$count = 54270;
	#10 counter$count = 54271;
	#10 counter$count = 54272;
	#10 counter$count = 54273;
	#10 counter$count = 54274;
	#10 counter$count = 54275;
	#10 counter$count = 54276;
	#10 counter$count = 54277;
	#10 counter$count = 54278;
	#10 counter$count = 54279;
	#10 counter$count = 54280;
	#10 counter$count = 54281;
	#10 counter$count = 54282;
	#10 counter$count = 54283;
	#10 counter$count = 54284;
	#10 counter$count = 54285;
	#10 counter$count = 54286;
	#10 counter$count = 54287;
	#10 counter$count = 54288;
	#10 counter$count = 54289;
	#10 counter$count = 54290;
	#10 counter$count = 54291;
	#10 counter$count = 54292;
	#10 counter$count = 54293;
	#10 counter$count = 54294;
	#10 counter$count = 54295;
	#10 counter$count = 54296;
	#10 counter$count = 54297;
	#10 counter$count = 54298;
	#10 counter$count = 54299;
	#10 counter$count = 54300;
	#10 counter$count = 54301;
	#10 counter$count = 54302;
	#10 counter$count = 54303;
	#10 counter$count = 54304;
	#10 counter$count = 54305;
	#10 counter$count = 54306;
	#10 counter$count = 54307;
	#10 counter$count = 54308;
	#10 counter$count = 54309;
	#10 counter$count = 54310;
	#10 counter$count = 54311;
	#10 counter$count = 54312;
	#10 counter$count = 54313;
	#10 counter$count = 54314;
	#10 counter$count = 54315;
	#10 counter$count = 54316;
	#10 counter$count = 54317;
	#10 counter$count = 54318;
	#10 counter$count = 54319;
	#10 counter$count = 54320;
	#10 counter$count = 54321;
	#10 counter$count = 54322;
	#10 counter$count = 54323;
	#10 counter$count = 54324;
	#10 counter$count = 54325;
	#10 counter$count = 54326;
	#10 counter$count = 54327;
	#10 counter$count = 54328;
	#10 counter$count = 54329;
	#10 counter$count = 54330;
	#10 counter$count = 54331;
	#10 counter$count = 54332;
	#10 counter$count = 54333;
	#10 counter$count = 54334;
	#10 counter$count = 54335;
	#10 counter$count = 54336;
	#10 counter$count = 54337;
	#10 counter$count = 54338;
	#10 counter$count = 54339;
	#10 counter$count = 54340;
	#10 counter$count = 54341;
	#10 counter$count = 54342;
	#10 counter$count = 54343;
	#10 counter$count = 54344;
	#10 counter$count = 54345;
	#10 counter$count = 54346;
	#10 counter$count = 54347;
	#10 counter$count = 54348;
	#10 counter$count = 54349;
	#10 counter$count = 54350;
	#10 counter$count = 54351;
	#10 counter$count = 54352;
	#10 counter$count = 54353;
	#10 counter$count = 54354;
	#10 counter$count = 54355;
	#10 counter$count = 54356;
	#10 counter$count = 54357;
	#10 counter$count = 54358;
	#10 counter$count = 54359;
	#10 counter$count = 54360;
	#10 counter$count = 54361;
	#10 counter$count = 54362;
	#10 counter$count = 54363;
	#10 counter$count = 54364;
	#10 counter$count = 54365;
	#10 counter$count = 54366;
	#10 counter$count = 54367;
	#10 counter$count = 54368;
	#10 counter$count = 54369;
	#10 counter$count = 54370;
	#10 counter$count = 54371;
	#10 counter$count = 54372;
	#10 counter$count = 54373;
	#10 counter$count = 54374;
	#10 counter$count = 54375;
	#10 counter$count = 54376;
	#10 counter$count = 54377;
	#10 counter$count = 54378;
	#10 counter$count = 54379;
	#10 counter$count = 54380;
	#10 counter$count = 54381;
	#10 counter$count = 54382;
	#10 counter$count = 54383;
	#10 counter$count = 54384;
	#10 counter$count = 54385;
	#10 counter$count = 54386;
	#10 counter$count = 54387;
	#10 counter$count = 54388;
	#10 counter$count = 54389;
	#10 counter$count = 54390;
	#10 counter$count = 54391;
	#10 counter$count = 54392;
	#10 counter$count = 54393;
	#10 counter$count = 54394;
	#10 counter$count = 54395;
	#10 counter$count = 54396;
	#10 counter$count = 54397;
	#10 counter$count = 54398;
	#10 counter$count = 54399;
	#10 counter$count = 54400;
	#10 counter$count = 54401;
	#10 counter$count = 54402;
	#10 counter$count = 54403;
	#10 counter$count = 54404;
	#10 counter$count = 54405;
	#10 counter$count = 54406;
	#10 counter$count = 54407;
	#10 counter$count = 54408;
	#10 counter$count = 54409;
	#10 counter$count = 54410;
	#10 counter$count = 54411;
	#10 counter$count = 54412;
	#10 counter$count = 54413;
	#10 counter$count = 54414;
	#10 counter$count = 54415;
	#10 counter$count = 54416;
	#10 counter$count = 54417;
	#10 counter$count = 54418;
	#10 counter$count = 54419;
	#10 counter$count = 54420;
	#10 counter$count = 54421;
	#10 counter$count = 54422;
	#10 counter$count = 54423;
	#10 counter$count = 54424;
	#10 counter$count = 54425;
	#10 counter$count = 54426;
	#10 counter$count = 54427;
	#10 counter$count = 54428;
	#10 counter$count = 54429;
	#10 counter$count = 54430;
	#10 counter$count = 54431;
	#10 counter$count = 54432;
	#10 counter$count = 54433;
	#10 counter$count = 54434;
	#10 counter$count = 54435;
	#10 counter$count = 54436;
	#10 counter$count = 54437;
	#10 counter$count = 54438;
	#10 counter$count = 54439;
	#10 counter$count = 54440;
	#10 counter$count = 54441;
	#10 counter$count = 54442;
	#10 counter$count = 54443;
	#10 counter$count = 54444;
	#10 counter$count = 54445;
	#10 counter$count = 54446;
	#10 counter$count = 54447;
	#10 counter$count = 54448;
	#10 counter$count = 54449;
	#10 counter$count = 54450;
	#10 counter$count = 54451;
	#10 counter$count = 54452;
	#10 counter$count = 54453;
	#10 counter$count = 54454;
	#10 counter$count = 54455;
	#10 counter$count = 54456;
	#10 counter$count = 54457;
	#10 counter$count = 54458;
	#10 counter$count = 54459;
	#10 counter$count = 54460;
	#10 counter$count = 54461;
	#10 counter$count = 54462;
	#10 counter$count = 54463;
	#10 counter$count = 54464;
	#10 counter$count = 54465;
	#10 counter$count = 54466;
	#10 counter$count = 54467;
	#10 counter$count = 54468;
	#10 counter$count = 54469;
	#10 counter$count = 54470;
	#10 counter$count = 54471;
	#10 counter$count = 54472;
	#10 counter$count = 54473;
	#10 counter$count = 54474;
	#10 counter$count = 54475;
	#10 counter$count = 54476;
	#10 counter$count = 54477;
	#10 counter$count = 54478;
	#10 counter$count = 54479;
	#10 counter$count = 54480;
	#10 counter$count = 54481;
	#10 counter$count = 54482;
	#10 counter$count = 54483;
	#10 counter$count = 54484;
	#10 counter$count = 54485;
	#10 counter$count = 54486;
	#10 counter$count = 54487;
	#10 counter$count = 54488;
	#10 counter$count = 54489;
	#10 counter$count = 54490;
	#10 counter$count = 54491;
	#10 counter$count = 54492;
	#10 counter$count = 54493;
	#10 counter$count = 54494;
	#10 counter$count = 54495;
	#10 counter$count = 54496;
	#10 counter$count = 54497;
	#10 counter$count = 54498;
	#10 counter$count = 54499;
	#10 counter$count = 54500;
	#10 counter$count = 54501;
	#10 counter$count = 54502;
	#10 counter$count = 54503;
	#10 counter$count = 54504;
	#10 counter$count = 54505;
	#10 counter$count = 54506;
	#10 counter$count = 54507;
	#10 counter$count = 54508;
	#10 counter$count = 54509;
	#10 counter$count = 54510;
	#10 counter$count = 54511;
	#10 counter$count = 54512;
	#10 counter$count = 54513;
	#10 counter$count = 54514;
	#10 counter$count = 54515;
	#10 counter$count = 54516;
	#10 counter$count = 54517;
	#10 counter$count = 54518;
	#10 counter$count = 54519;
	#10 counter$count = 54520;
	#10 counter$count = 54521;
	#10 counter$count = 54522;
	#10 counter$count = 54523;
	#10 counter$count = 54524;
	#10 counter$count = 54525;
	#10 counter$count = 54526;
	#10 counter$count = 54527;
	#10 counter$count = 54528;
	#10 counter$count = 54529;
	#10 counter$count = 54530;
	#10 counter$count = 54531;
	#10 counter$count = 54532;
	#10 counter$count = 54533;
	#10 counter$count = 54534;
	#10 counter$count = 54535;
	#10 counter$count = 54536;
	#10 counter$count = 54537;
	#10 counter$count = 54538;
	#10 counter$count = 54539;
	#10 counter$count = 54540;
	#10 counter$count = 54541;
	#10 counter$count = 54542;
	#10 counter$count = 54543;
	#10 counter$count = 54544;
	#10 counter$count = 54545;
	#10 counter$count = 54546;
	#10 counter$count = 54547;
	#10 counter$count = 54548;
	#10 counter$count = 54549;
	#10 counter$count = 54550;
	#10 counter$count = 54551;
	#10 counter$count = 54552;
	#10 counter$count = 54553;
	#10 counter$count = 54554;
	#10 counter$count = 54555;
	#10 counter$count = 54556;
	#10 counter$count = 54557;
	#10 counter$count = 54558;
	#10 counter$count = 54559;
	#10 counter$count = 54560;
	#10 counter$count = 54561;
	#10 counter$count = 54562;
	#10 counter$count = 54563;
	#10 counter$count = 54564;
	#10 counter$count = 54565;
	#10 counter$count = 54566;
	#10 counter$count = 54567;
	#10 counter$count = 54568;
	#10 counter$count = 54569;
	#10 counter$count = 54570;
	#10 counter$count = 54571;
	#10 counter$count = 54572;
	#10 counter$count = 54573;
	#10 counter$count = 54574;
	#10 counter$count = 54575;
	#10 counter$count = 54576;
	#10 counter$count = 54577;
	#10 counter$count = 54578;
	#10 counter$count = 54579;
	#10 counter$count = 54580;
	#10 counter$count = 54581;
	#10 counter$count = 54582;
	#10 counter$count = 54583;
	#10 counter$count = 54584;
	#10 counter$count = 54585;
	#10 counter$count = 54586;
	#10 counter$count = 54587;
	#10 counter$count = 54588;
	#10 counter$count = 54589;
	#10 counter$count = 54590;
	#10 counter$count = 54591;
	#10 counter$count = 54592;
	#10 counter$count = 54593;
	#10 counter$count = 54594;
	#10 counter$count = 54595;
	#10 counter$count = 54596;
	#10 counter$count = 54597;
	#10 counter$count = 54598;
	#10 counter$count = 54599;
	#10 counter$count = 54600;
	#10 counter$count = 54601;
	#10 counter$count = 54602;
	#10 counter$count = 54603;
	#10 counter$count = 54604;
	#10 counter$count = 54605;
	#10 counter$count = 54606;
	#10 counter$count = 54607;
	#10 counter$count = 54608;
	#10 counter$count = 54609;
	#10 counter$count = 54610;
	#10 counter$count = 54611;
	#10 counter$count = 54612;
	#10 counter$count = 54613;
	#10 counter$count = 54614;
	#10 counter$count = 54615;
	#10 counter$count = 54616;
	#10 counter$count = 54617;
	#10 counter$count = 54618;
	#10 counter$count = 54619;
	#10 counter$count = 54620;
	#10 counter$count = 54621;
	#10 counter$count = 54622;
	#10 counter$count = 54623;
	#10 counter$count = 54624;
	#10 counter$count = 54625;
	#10 counter$count = 54626;
	#10 counter$count = 54627;
	#10 counter$count = 54628;
	#10 counter$count = 54629;
	#10 counter$count = 54630;
	#10 counter$count = 54631;
	#10 counter$count = 54632;
	#10 counter$count = 54633;
	#10 counter$count = 54634;
	#10 counter$count = 54635;
	#10 counter$count = 54636;
	#10 counter$count = 54637;
	#10 counter$count = 54638;
	#10 counter$count = 54639;
	#10 counter$count = 54640;
	#10 counter$count = 54641;
	#10 counter$count = 54642;
	#10 counter$count = 54643;
	#10 counter$count = 54644;
	#10 counter$count = 54645;
	#10 counter$count = 54646;
	#10 counter$count = 54647;
	#10 counter$count = 54648;
	#10 counter$count = 54649;
	#10 counter$count = 54650;
	#10 counter$count = 54651;
	#10 counter$count = 54652;
	#10 counter$count = 54653;
	#10 counter$count = 54654;
	#10 counter$count = 54655;
	#10 counter$count = 54656;
	#10 counter$count = 54657;
	#10 counter$count = 54658;
	#10 counter$count = 54659;
	#10 counter$count = 54660;
	#10 counter$count = 54661;
	#10 counter$count = 54662;
	#10 counter$count = 54663;
	#10 counter$count = 54664;
	#10 counter$count = 54665;
	#10 counter$count = 54666;
	#10 counter$count = 54667;
	#10 counter$count = 54668;
	#10 counter$count = 54669;
	#10 counter$count = 54670;
	#10 counter$count = 54671;
	#10 counter$count = 54672;
	#10 counter$count = 54673;
	#10 counter$count = 54674;
	#10 counter$count = 54675;
	#10 counter$count = 54676;
	#10 counter$count = 54677;
	#10 counter$count = 54678;
	#10 counter$count = 54679;
	#10 counter$count = 54680;
	#10 counter$count = 54681;
	#10 counter$count = 54682;
	#10 counter$count = 54683;
	#10 counter$count = 54684;
	#10 counter$count = 54685;
	#10 counter$count = 54686;
	#10 counter$count = 54687;
	#10 counter$count = 54688;
	#10 counter$count = 54689;
	#10 counter$count = 54690;
	#10 counter$count = 54691;
	#10 counter$count = 54692;
	#10 counter$count = 54693;
	#10 counter$count = 54694;
	#10 counter$count = 54695;
	#10 counter$count = 54696;
	#10 counter$count = 54697;
	#10 counter$count = 54698;
	#10 counter$count = 54699;
	#10 counter$count = 54700;
	#10 counter$count = 54701;
	#10 counter$count = 54702;
	#10 counter$count = 54703;
	#10 counter$count = 54704;
	#10 counter$count = 54705;
	#10 counter$count = 54706;
	#10 counter$count = 54707;
	#10 counter$count = 54708;
	#10 counter$count = 54709;
	#10 counter$count = 54710;
	#10 counter$count = 54711;
	#10 counter$count = 54712;
	#10 counter$count = 54713;
	#10 counter$count = 54714;
	#10 counter$count = 54715;
	#10 counter$count = 54716;
	#10 counter$count = 54717;
	#10 counter$count = 54718;
	#10 counter$count = 54719;
	#10 counter$count = 54720;
	#10 counter$count = 54721;
	#10 counter$count = 54722;
	#10 counter$count = 54723;
	#10 counter$count = 54724;
	#10 counter$count = 54725;
	#10 counter$count = 54726;
	#10 counter$count = 54727;
	#10 counter$count = 54728;
	#10 counter$count = 54729;
	#10 counter$count = 54730;
	#10 counter$count = 54731;
	#10 counter$count = 54732;
	#10 counter$count = 54733;
	#10 counter$count = 54734;
	#10 counter$count = 54735;
	#10 counter$count = 54736;
	#10 counter$count = 54737;
	#10 counter$count = 54738;
	#10 counter$count = 54739;
	#10 counter$count = 54740;
	#10 counter$count = 54741;
	#10 counter$count = 54742;
	#10 counter$count = 54743;
	#10 counter$count = 54744;
	#10 counter$count = 54745;
	#10 counter$count = 54746;
	#10 counter$count = 54747;
	#10 counter$count = 54748;
	#10 counter$count = 54749;
	#10 counter$count = 54750;
	#10 counter$count = 54751;
	#10 counter$count = 54752;
	#10 counter$count = 54753;
	#10 counter$count = 54754;
	#10 counter$count = 54755;
	#10 counter$count = 54756;
	#10 counter$count = 54757;
	#10 counter$count = 54758;
	#10 counter$count = 54759;
	#10 counter$count = 54760;
	#10 counter$count = 54761;
	#10 counter$count = 54762;
	#10 counter$count = 54763;
	#10 counter$count = 54764;
	#10 counter$count = 54765;
	#10 counter$count = 54766;
	#10 counter$count = 54767;
	#10 counter$count = 54768;
	#10 counter$count = 54769;
	#10 counter$count = 54770;
	#10 counter$count = 54771;
	#10 counter$count = 54772;
	#10 counter$count = 54773;
	#10 counter$count = 54774;
	#10 counter$count = 54775;
	#10 counter$count = 54776;
	#10 counter$count = 54777;
	#10 counter$count = 54778;
	#10 counter$count = 54779;
	#10 counter$count = 54780;
	#10 counter$count = 54781;
	#10 counter$count = 54782;
	#10 counter$count = 54783;
	#10 counter$count = 54784;
	#10 counter$count = 54785;
	#10 counter$count = 54786;
	#10 counter$count = 54787;
	#10 counter$count = 54788;
	#10 counter$count = 54789;
	#10 counter$count = 54790;
	#10 counter$count = 54791;
	#10 counter$count = 54792;
	#10 counter$count = 54793;
	#10 counter$count = 54794;
	#10 counter$count = 54795;
	#10 counter$count = 54796;
	#10 counter$count = 54797;
	#10 counter$count = 54798;
	#10 counter$count = 54799;
	#10 counter$count = 54800;
	#10 counter$count = 54801;
	#10 counter$count = 54802;
	#10 counter$count = 54803;
	#10 counter$count = 54804;
	#10 counter$count = 54805;
	#10 counter$count = 54806;
	#10 counter$count = 54807;
	#10 counter$count = 54808;
	#10 counter$count = 54809;
	#10 counter$count = 54810;
	#10 counter$count = 54811;
	#10 counter$count = 54812;
	#10 counter$count = 54813;
	#10 counter$count = 54814;
	#10 counter$count = 54815;
	#10 counter$count = 54816;
	#10 counter$count = 54817;
	#10 counter$count = 54818;
	#10 counter$count = 54819;
	#10 counter$count = 54820;
	#10 counter$count = 54821;
	#10 counter$count = 54822;
	#10 counter$count = 54823;
	#10 counter$count = 54824;
	#10 counter$count = 54825;
	#10 counter$count = 54826;
	#10 counter$count = 54827;
	#10 counter$count = 54828;
	#10 counter$count = 54829;
	#10 counter$count = 54830;
	#10 counter$count = 54831;
	#10 counter$count = 54832;
	#10 counter$count = 54833;
	#10 counter$count = 54834;
	#10 counter$count = 54835;
	#10 counter$count = 54836;
	#10 counter$count = 54837;
	#10 counter$count = 54838;
	#10 counter$count = 54839;
	#10 counter$count = 54840;
	#10 counter$count = 54841;
	#10 counter$count = 54842;
	#10 counter$count = 54843;
	#10 counter$count = 54844;
	#10 counter$count = 54845;
	#10 counter$count = 54846;
	#10 counter$count = 54847;
	#10 counter$count = 54848;
	#10 counter$count = 54849;
	#10 counter$count = 54850;
	#10 counter$count = 54851;
	#10 counter$count = 54852;
	#10 counter$count = 54853;
	#10 counter$count = 54854;
	#10 counter$count = 54855;
	#10 counter$count = 54856;
	#10 counter$count = 54857;
	#10 counter$count = 54858;
	#10 counter$count = 54859;
	#10 counter$count = 54860;
	#10 counter$count = 54861;
	#10 counter$count = 54862;
	#10 counter$count = 54863;
	#10 counter$count = 54864;
	#10 counter$count = 54865;
	#10 counter$count = 54866;
	#10 counter$count = 54867;
	#10 counter$count = 54868;
	#10 counter$count = 54869;
	#10 counter$count = 54870;
	#10 counter$count = 54871;
	#10 counter$count = 54872;
	#10 counter$count = 54873;
	#10 counter$count = 54874;
	#10 counter$count = 54875;
	#10 counter$count = 54876;
	#10 counter$count = 54877;
	#10 counter$count = 54878;
	#10 counter$count = 54879;
	#10 counter$count = 54880;
	#10 counter$count = 54881;
	#10 counter$count = 54882;
	#10 counter$count = 54883;
	#10 counter$count = 54884;
	#10 counter$count = 54885;
	#10 counter$count = 54886;
	#10 counter$count = 54887;
	#10 counter$count = 54888;
	#10 counter$count = 54889;
	#10 counter$count = 54890;
	#10 counter$count = 54891;
	#10 counter$count = 54892;
	#10 counter$count = 54893;
	#10 counter$count = 54894;
	#10 counter$count = 54895;
	#10 counter$count = 54896;
	#10 counter$count = 54897;
	#10 counter$count = 54898;
	#10 counter$count = 54899;
	#10 counter$count = 54900;
	#10 counter$count = 54901;
	#10 counter$count = 54902;
	#10 counter$count = 54903;
	#10 counter$count = 54904;
	#10 counter$count = 54905;
	#10 counter$count = 54906;
	#10 counter$count = 54907;
	#10 counter$count = 54908;
	#10 counter$count = 54909;
	#10 counter$count = 54910;
	#10 counter$count = 54911;
	#10 counter$count = 54912;
	#10 counter$count = 54913;
	#10 counter$count = 54914;
	#10 counter$count = 54915;
	#10 counter$count = 54916;
	#10 counter$count = 54917;
	#10 counter$count = 54918;
	#10 counter$count = 54919;
	#10 counter$count = 54920;
	#10 counter$count = 54921;
	#10 counter$count = 54922;
	#10 counter$count = 54923;
	#10 counter$count = 54924;
	#10 counter$count = 54925;
	#10 counter$count = 54926;
	#10 counter$count = 54927;
	#10 counter$count = 54928;
	#10 counter$count = 54929;
	#10 counter$count = 54930;
	#10 counter$count = 54931;
	#10 counter$count = 54932;
	#10 counter$count = 54933;
	#10 counter$count = 54934;
	#10 counter$count = 54935;
	#10 counter$count = 54936;
	#10 counter$count = 54937;
	#10 counter$count = 54938;
	#10 counter$count = 54939;
	#10 counter$count = 54940;
	#10 counter$count = 54941;
	#10 counter$count = 54942;
	#10 counter$count = 54943;
	#10 counter$count = 54944;
	#10 counter$count = 54945;
	#10 counter$count = 54946;
	#10 counter$count = 54947;
	#10 counter$count = 54948;
	#10 counter$count = 54949;
	#10 counter$count = 54950;
	#10 counter$count = 54951;
	#10 counter$count = 54952;
	#10 counter$count = 54953;
	#10 counter$count = 54954;
	#10 counter$count = 54955;
	#10 counter$count = 54956;
	#10 counter$count = 54957;
	#10 counter$count = 54958;
	#10 counter$count = 54959;
	#10 counter$count = 54960;
	#10 counter$count = 54961;
	#10 counter$count = 54962;
	#10 counter$count = 54963;
	#10 counter$count = 54964;
	#10 counter$count = 54965;
	#10 counter$count = 54966;
	#10 counter$count = 54967;
	#10 counter$count = 54968;
	#10 counter$count = 54969;
	#10 counter$count = 54970;
	#10 counter$count = 54971;
	#10 counter$count = 54972;
	#10 counter$count = 54973;
	#10 counter$count = 54974;
	#10 counter$count = 54975;
	#10 counter$count = 54976;
	#10 counter$count = 54977;
	#10 counter$count = 54978;
	#10 counter$count = 54979;
	#10 counter$count = 54980;
	#10 counter$count = 54981;
	#10 counter$count = 54982;
	#10 counter$count = 54983;
	#10 counter$count = 54984;
	#10 counter$count = 54985;
	#10 counter$count = 54986;
	#10 counter$count = 54987;
	#10 counter$count = 54988;
	#10 counter$count = 54989;
	#10 counter$count = 54990;
	#10 counter$count = 54991;
	#10 counter$count = 54992;
	#10 counter$count = 54993;
	#10 counter$count = 54994;
	#10 counter$count = 54995;
	#10 counter$count = 54996;
	#10 counter$count = 54997;
	#10 counter$count = 54998;
	#10 counter$count = 54999;
	#10 counter$count = 55000;
	#10 counter$count = 55001;
	#10 counter$count = 55002;
	#10 counter$count = 55003;
	#10 counter$count = 55004;
	#10 counter$count = 55005;
	#10 counter$count = 55006;
	#10 counter$count = 55007;
	#10 counter$count = 55008;
	#10 counter$count = 55009;
	#10 counter$count = 55010;
	#10 counter$count = 55011;
	#10 counter$count = 55012;
	#10 counter$count = 55013;
	#10 counter$count = 55014;
	#10 counter$count = 55015;
	#10 counter$count = 55016;
	#10 counter$count = 55017;
	#10 counter$count = 55018;
	#10 counter$count = 55019;
	#10 counter$count = 55020;
	#10 counter$count = 55021;
	#10 counter$count = 55022;
	#10 counter$count = 55023;
	#10 counter$count = 55024;
	#10 counter$count = 55025;
	#10 counter$count = 55026;
	#10 counter$count = 55027;
	#10 counter$count = 55028;
	#10 counter$count = 55029;
	#10 counter$count = 55030;
	#10 counter$count = 55031;
	#10 counter$count = 55032;
	#10 counter$count = 55033;
	#10 counter$count = 55034;
	#10 counter$count = 55035;
	#10 counter$count = 55036;
	#10 counter$count = 55037;
	#10 counter$count = 55038;
	#10 counter$count = 55039;
	#10 counter$count = 55040;
	#10 counter$count = 55041;
	#10 counter$count = 55042;
	#10 counter$count = 55043;
	#10 counter$count = 55044;
	#10 counter$count = 55045;
	#10 counter$count = 55046;
	#10 counter$count = 55047;
	#10 counter$count = 55048;
	#10 counter$count = 55049;
	#10 counter$count = 55050;
	#10 counter$count = 55051;
	#10 counter$count = 55052;
	#10 counter$count = 55053;
	#10 counter$count = 55054;
	#10 counter$count = 55055;
	#10 counter$count = 55056;
	#10 counter$count = 55057;
	#10 counter$count = 55058;
	#10 counter$count = 55059;
	#10 counter$count = 55060;
	#10 counter$count = 55061;
	#10 counter$count = 55062;
	#10 counter$count = 55063;
	#10 counter$count = 55064;
	#10 counter$count = 55065;
	#10 counter$count = 55066;
	#10 counter$count = 55067;
	#10 counter$count = 55068;
	#10 counter$count = 55069;
	#10 counter$count = 55070;
	#10 counter$count = 55071;
	#10 counter$count = 55072;
	#10 counter$count = 55073;
	#10 counter$count = 55074;
	#10 counter$count = 55075;
	#10 counter$count = 55076;
	#10 counter$count = 55077;
	#10 counter$count = 55078;
	#10 counter$count = 55079;
	#10 counter$count = 55080;
	#10 counter$count = 55081;
	#10 counter$count = 55082;
	#10 counter$count = 55083;
	#10 counter$count = 55084;
	#10 counter$count = 55085;
	#10 counter$count = 55086;
	#10 counter$count = 55087;
	#10 counter$count = 55088;
	#10 counter$count = 55089;
	#10 counter$count = 55090;
	#10 counter$count = 55091;
	#10 counter$count = 55092;
	#10 counter$count = 55093;
	#10 counter$count = 55094;
	#10 counter$count = 55095;
	#10 counter$count = 55096;
	#10 counter$count = 55097;
	#10 counter$count = 55098;
	#10 counter$count = 55099;
	#10 counter$count = 55100;
	#10 counter$count = 55101;
	#10 counter$count = 55102;
	#10 counter$count = 55103;
	#10 counter$count = 55104;
	#10 counter$count = 55105;
	#10 counter$count = 55106;
	#10 counter$count = 55107;
	#10 counter$count = 55108;
	#10 counter$count = 55109;
	#10 counter$count = 55110;
	#10 counter$count = 55111;
	#10 counter$count = 55112;
	#10 counter$count = 55113;
	#10 counter$count = 55114;
	#10 counter$count = 55115;
	#10 counter$count = 55116;
	#10 counter$count = 55117;
	#10 counter$count = 55118;
	#10 counter$count = 55119;
	#10 counter$count = 55120;
	#10 counter$count = 55121;
	#10 counter$count = 55122;
	#10 counter$count = 55123;
	#10 counter$count = 55124;
	#10 counter$count = 55125;
	#10 counter$count = 55126;
	#10 counter$count = 55127;
	#10 counter$count = 55128;
	#10 counter$count = 55129;
	#10 counter$count = 55130;
	#10 counter$count = 55131;
	#10 counter$count = 55132;
	#10 counter$count = 55133;
	#10 counter$count = 55134;
	#10 counter$count = 55135;
	#10 counter$count = 55136;
	#10 counter$count = 55137;
	#10 counter$count = 55138;
	#10 counter$count = 55139;
	#10 counter$count = 55140;
	#10 counter$count = 55141;
	#10 counter$count = 55142;
	#10 counter$count = 55143;
	#10 counter$count = 55144;
	#10 counter$count = 55145;
	#10 counter$count = 55146;
	#10 counter$count = 55147;
	#10 counter$count = 55148;
	#10 counter$count = 55149;
	#10 counter$count = 55150;
	#10 counter$count = 55151;
	#10 counter$count = 55152;
	#10 counter$count = 55153;
	#10 counter$count = 55154;
	#10 counter$count = 55155;
	#10 counter$count = 55156;
	#10 counter$count = 55157;
	#10 counter$count = 55158;
	#10 counter$count = 55159;
	#10 counter$count = 55160;
	#10 counter$count = 55161;
	#10 counter$count = 55162;
	#10 counter$count = 55163;
	#10 counter$count = 55164;
	#10 counter$count = 55165;
	#10 counter$count = 55166;
	#10 counter$count = 55167;
	#10 counter$count = 55168;
	#10 counter$count = 55169;
	#10 counter$count = 55170;
	#10 counter$count = 55171;
	#10 counter$count = 55172;
	#10 counter$count = 55173;
	#10 counter$count = 55174;
	#10 counter$count = 55175;
	#10 counter$count = 55176;
	#10 counter$count = 55177;
	#10 counter$count = 55178;
	#10 counter$count = 55179;
	#10 counter$count = 55180;
	#10 counter$count = 55181;
	#10 counter$count = 55182;
	#10 counter$count = 55183;
	#10 counter$count = 55184;
	#10 counter$count = 55185;
	#10 counter$count = 55186;
	#10 counter$count = 55187;
	#10 counter$count = 55188;
	#10 counter$count = 55189;
	#10 counter$count = 55190;
	#10 counter$count = 55191;
	#10 counter$count = 55192;
	#10 counter$count = 55193;
	#10 counter$count = 55194;
	#10 counter$count = 55195;
	#10 counter$count = 55196;
	#10 counter$count = 55197;
	#10 counter$count = 55198;
	#10 counter$count = 55199;
	#10 counter$count = 55200;
	#10 counter$count = 55201;
	#10 counter$count = 55202;
	#10 counter$count = 55203;
	#10 counter$count = 55204;
	#10 counter$count = 55205;
	#10 counter$count = 55206;
	#10 counter$count = 55207;
	#10 counter$count = 55208;
	#10 counter$count = 55209;
	#10 counter$count = 55210;
	#10 counter$count = 55211;
	#10 counter$count = 55212;
	#10 counter$count = 55213;
	#10 counter$count = 55214;
	#10 counter$count = 55215;
	#10 counter$count = 55216;
	#10 counter$count = 55217;
	#10 counter$count = 55218;
	#10 counter$count = 55219;
	#10 counter$count = 55220;
	#10 counter$count = 55221;
	#10 counter$count = 55222;
	#10 counter$count = 55223;
	#10 counter$count = 55224;
	#10 counter$count = 55225;
	#10 counter$count = 55226;
	#10 counter$count = 55227;
	#10 counter$count = 55228;
	#10 counter$count = 55229;
	#10 counter$count = 55230;
	#10 counter$count = 55231;
	#10 counter$count = 55232;
	#10 counter$count = 55233;
	#10 counter$count = 55234;
	#10 counter$count = 55235;
	#10 counter$count = 55236;
	#10 counter$count = 55237;
	#10 counter$count = 55238;
	#10 counter$count = 55239;
	#10 counter$count = 55240;
	#10 counter$count = 55241;
	#10 counter$count = 55242;
	#10 counter$count = 55243;
	#10 counter$count = 55244;
	#10 counter$count = 55245;
	#10 counter$count = 55246;
	#10 counter$count = 55247;
	#10 counter$count = 55248;
	#10 counter$count = 55249;
	#10 counter$count = 55250;
	#10 counter$count = 55251;
	#10 counter$count = 55252;
	#10 counter$count = 55253;
	#10 counter$count = 55254;
	#10 counter$count = 55255;
	#10 counter$count = 55256;
	#10 counter$count = 55257;
	#10 counter$count = 55258;
	#10 counter$count = 55259;
	#10 counter$count = 55260;
	#10 counter$count = 55261;
	#10 counter$count = 55262;
	#10 counter$count = 55263;
	#10 counter$count = 55264;
	#10 counter$count = 55265;
	#10 counter$count = 55266;
	#10 counter$count = 55267;
	#10 counter$count = 55268;
	#10 counter$count = 55269;
	#10 counter$count = 55270;
	#10 counter$count = 55271;
	#10 counter$count = 55272;
	#10 counter$count = 55273;
	#10 counter$count = 55274;
	#10 counter$count = 55275;
	#10 counter$count = 55276;
	#10 counter$count = 55277;
	#10 counter$count = 55278;
	#10 counter$count = 55279;
	#10 counter$count = 55280;
	#10 counter$count = 55281;
	#10 counter$count = 55282;
	#10 counter$count = 55283;
	#10 counter$count = 55284;
	#10 counter$count = 55285;
	#10 counter$count = 55286;
	#10 counter$count = 55287;
	#10 counter$count = 55288;
	#10 counter$count = 55289;
	#10 counter$count = 55290;
	#10 counter$count = 55291;
	#10 counter$count = 55292;
	#10 counter$count = 55293;
	#10 counter$count = 55294;
	#10 counter$count = 55295;
	#10 counter$count = 55296;
	#10 counter$count = 55297;
	#10 counter$count = 55298;
	#10 counter$count = 55299;
	#10 counter$count = 55300;
	#10 counter$count = 55301;
	#10 counter$count = 55302;
	#10 counter$count = 55303;
	#10 counter$count = 55304;
	#10 counter$count = 55305;
	#10 counter$count = 55306;
	#10 counter$count = 55307;
	#10 counter$count = 55308;
	#10 counter$count = 55309;
	#10 counter$count = 55310;
	#10 counter$count = 55311;
	#10 counter$count = 55312;
	#10 counter$count = 55313;
	#10 counter$count = 55314;
	#10 counter$count = 55315;
	#10 counter$count = 55316;
	#10 counter$count = 55317;
	#10 counter$count = 55318;
	#10 counter$count = 55319;
	#10 counter$count = 55320;
	#10 counter$count = 55321;
	#10 counter$count = 55322;
	#10 counter$count = 55323;
	#10 counter$count = 55324;
	#10 counter$count = 55325;
	#10 counter$count = 55326;
	#10 counter$count = 55327;
	#10 counter$count = 55328;
	#10 counter$count = 55329;
	#10 counter$count = 55330;
	#10 counter$count = 55331;
	#10 counter$count = 55332;
	#10 counter$count = 55333;
	#10 counter$count = 55334;
	#10 counter$count = 55335;
	#10 counter$count = 55336;
	#10 counter$count = 55337;
	#10 counter$count = 55338;
	#10 counter$count = 55339;
	#10 counter$count = 55340;
	#10 counter$count = 55341;
	#10 counter$count = 55342;
	#10 counter$count = 55343;
	#10 counter$count = 55344;
	#10 counter$count = 55345;
	#10 counter$count = 55346;
	#10 counter$count = 55347;
	#10 counter$count = 55348;
	#10 counter$count = 55349;
	#10 counter$count = 55350;
	#10 counter$count = 55351;
	#10 counter$count = 55352;
	#10 counter$count = 55353;
	#10 counter$count = 55354;
	#10 counter$count = 55355;
	#10 counter$count = 55356;
	#10 counter$count = 55357;
	#10 counter$count = 55358;
	#10 counter$count = 55359;
	#10 counter$count = 55360;
	#10 counter$count = 55361;
	#10 counter$count = 55362;
	#10 counter$count = 55363;
	#10 counter$count = 55364;
	#10 counter$count = 55365;
	#10 counter$count = 55366;
	#10 counter$count = 55367;
	#10 counter$count = 55368;
	#10 counter$count = 55369;
	#10 counter$count = 55370;
	#10 counter$count = 55371;
	#10 counter$count = 55372;
	#10 counter$count = 55373;
	#10 counter$count = 55374;
	#10 counter$count = 55375;
	#10 counter$count = 55376;
	#10 counter$count = 55377;
	#10 counter$count = 55378;
	#10 counter$count = 55379;
	#10 counter$count = 55380;
	#10 counter$count = 55381;
	#10 counter$count = 55382;
	#10 counter$count = 55383;
	#10 counter$count = 55384;
	#10 counter$count = 55385;
	#10 counter$count = 55386;
	#10 counter$count = 55387;
	#10 counter$count = 55388;
	#10 counter$count = 55389;
	#10 counter$count = 55390;
	#10 counter$count = 55391;
	#10 counter$count = 55392;
	#10 counter$count = 55393;
	#10 counter$count = 55394;
	#10 counter$count = 55395;
	#10 counter$count = 55396;
	#10 counter$count = 55397;
	#10 counter$count = 55398;
	#10 counter$count = 55399;
	#10 counter$count = 55400;
	#10 counter$count = 55401;
	#10 counter$count = 55402;
	#10 counter$count = 55403;
	#10 counter$count = 55404;
	#10 counter$count = 55405;
	#10 counter$count = 55406;
	#10 counter$count = 55407;
	#10 counter$count = 55408;
	#10 counter$count = 55409;
	#10 counter$count = 55410;
	#10 counter$count = 55411;
	#10 counter$count = 55412;
	#10 counter$count = 55413;
	#10 counter$count = 55414;
	#10 counter$count = 55415;
	#10 counter$count = 55416;
	#10 counter$count = 55417;
	#10 counter$count = 55418;
	#10 counter$count = 55419;
	#10 counter$count = 55420;
	#10 counter$count = 55421;
	#10 counter$count = 55422;
	#10 counter$count = 55423;
	#10 counter$count = 55424;
	#10 counter$count = 55425;
	#10 counter$count = 55426;
	#10 counter$count = 55427;
	#10 counter$count = 55428;
	#10 counter$count = 55429;
	#10 counter$count = 55430;
	#10 counter$count = 55431;
	#10 counter$count = 55432;
	#10 counter$count = 55433;
	#10 counter$count = 55434;
	#10 counter$count = 55435;
	#10 counter$count = 55436;
	#10 counter$count = 55437;
	#10 counter$count = 55438;
	#10 counter$count = 55439;
	#10 counter$count = 55440;
	#10 counter$count = 55441;
	#10 counter$count = 55442;
	#10 counter$count = 55443;
	#10 counter$count = 55444;
	#10 counter$count = 55445;
	#10 counter$count = 55446;
	#10 counter$count = 55447;
	#10 counter$count = 55448;
	#10 counter$count = 55449;
	#10 counter$count = 55450;
	#10 counter$count = 55451;
	#10 counter$count = 55452;
	#10 counter$count = 55453;
	#10 counter$count = 55454;
	#10 counter$count = 55455;
	#10 counter$count = 55456;
	#10 counter$count = 55457;
	#10 counter$count = 55458;
	#10 counter$count = 55459;
	#10 counter$count = 55460;
	#10 counter$count = 55461;
	#10 counter$count = 55462;
	#10 counter$count = 55463;
	#10 counter$count = 55464;
	#10 counter$count = 55465;
	#10 counter$count = 55466;
	#10 counter$count = 55467;
	#10 counter$count = 55468;
	#10 counter$count = 55469;
	#10 counter$count = 55470;
	#10 counter$count = 55471;
	#10 counter$count = 55472;
	#10 counter$count = 55473;
	#10 counter$count = 55474;
	#10 counter$count = 55475;
	#10 counter$count = 55476;
	#10 counter$count = 55477;
	#10 counter$count = 55478;
	#10 counter$count = 55479;
	#10 counter$count = 55480;
	#10 counter$count = 55481;
	#10 counter$count = 55482;
	#10 counter$count = 55483;
	#10 counter$count = 55484;
	#10 counter$count = 55485;
	#10 counter$count = 55486;
	#10 counter$count = 55487;
	#10 counter$count = 55488;
	#10 counter$count = 55489;
	#10 counter$count = 55490;
	#10 counter$count = 55491;
	#10 counter$count = 55492;
	#10 counter$count = 55493;
	#10 counter$count = 55494;
	#10 counter$count = 55495;
	#10 counter$count = 55496;
	#10 counter$count = 55497;
	#10 counter$count = 55498;
	#10 counter$count = 55499;
	#10 counter$count = 55500;
	#10 counter$count = 55501;
	#10 counter$count = 55502;
	#10 counter$count = 55503;
	#10 counter$count = 55504;
	#10 counter$count = 55505;
	#10 counter$count = 55506;
	#10 counter$count = 55507;
	#10 counter$count = 55508;
	#10 counter$count = 55509;
	#10 counter$count = 55510;
	#10 counter$count = 55511;
	#10 counter$count = 55512;
	#10 counter$count = 55513;
	#10 counter$count = 55514;
	#10 counter$count = 55515;
	#10 counter$count = 55516;
	#10 counter$count = 55517;
	#10 counter$count = 55518;
	#10 counter$count = 55519;
	#10 counter$count = 55520;
	#10 counter$count = 55521;
	#10 counter$count = 55522;
	#10 counter$count = 55523;
	#10 counter$count = 55524;
	#10 counter$count = 55525;
	#10 counter$count = 55526;
	#10 counter$count = 55527;
	#10 counter$count = 55528;
	#10 counter$count = 55529;
	#10 counter$count = 55530;
	#10 counter$count = 55531;
	#10 counter$count = 55532;
	#10 counter$count = 55533;
	#10 counter$count = 55534;
	#10 counter$count = 55535;
	#10 counter$count = 55536;
	#10 counter$count = 55537;
	#10 counter$count = 55538;
	#10 counter$count = 55539;
	#10 counter$count = 55540;
	#10 counter$count = 55541;
	#10 counter$count = 55542;
	#10 counter$count = 55543;
	#10 counter$count = 55544;
	#10 counter$count = 55545;
	#10 counter$count = 55546;
	#10 counter$count = 55547;
	#10 counter$count = 55548;
	#10 counter$count = 55549;
	#10 counter$count = 55550;
	#10 counter$count = 55551;
	#10 counter$count = 55552;
	#10 counter$count = 55553;
	#10 counter$count = 55554;
	#10 counter$count = 55555;
	#10 counter$count = 55556;
	#10 counter$count = 55557;
	#10 counter$count = 55558;
	#10 counter$count = 55559;
	#10 counter$count = 55560;
	#10 counter$count = 55561;
	#10 counter$count = 55562;
	#10 counter$count = 55563;
	#10 counter$count = 55564;
	#10 counter$count = 55565;
	#10 counter$count = 55566;
	#10 counter$count = 55567;
	#10 counter$count = 55568;
	#10 counter$count = 55569;
	#10 counter$count = 55570;
	#10 counter$count = 55571;
	#10 counter$count = 55572;
	#10 counter$count = 55573;
	#10 counter$count = 55574;
	#10 counter$count = 55575;
	#10 counter$count = 55576;
	#10 counter$count = 55577;
	#10 counter$count = 55578;
	#10 counter$count = 55579;
	#10 counter$count = 55580;
	#10 counter$count = 55581;
	#10 counter$count = 55582;
	#10 counter$count = 55583;
	#10 counter$count = 55584;
	#10 counter$count = 55585;
	#10 counter$count = 55586;
	#10 counter$count = 55587;
	#10 counter$count = 55588;
	#10 counter$count = 55589;
	#10 counter$count = 55590;
	#10 counter$count = 55591;
	#10 counter$count = 55592;
	#10 counter$count = 55593;
	#10 counter$count = 55594;
	#10 counter$count = 55595;
	#10 counter$count = 55596;
	#10 counter$count = 55597;
	#10 counter$count = 55598;
	#10 counter$count = 55599;
	#10 counter$count = 55600;
	#10 counter$count = 55601;
	#10 counter$count = 55602;
	#10 counter$count = 55603;
	#10 counter$count = 55604;
	#10 counter$count = 55605;
	#10 counter$count = 55606;
	#10 counter$count = 55607;
	#10 counter$count = 55608;
	#10 counter$count = 55609;
	#10 counter$count = 55610;
	#10 counter$count = 55611;
	#10 counter$count = 55612;
	#10 counter$count = 55613;
	#10 counter$count = 55614;
	#10 counter$count = 55615;
	#10 counter$count = 55616;
	#10 counter$count = 55617;
	#10 counter$count = 55618;
	#10 counter$count = 55619;
	#10 counter$count = 55620;
	#10 counter$count = 55621;
	#10 counter$count = 55622;
	#10 counter$count = 55623;
	#10 counter$count = 55624;
	#10 counter$count = 55625;
	#10 counter$count = 55626;
	#10 counter$count = 55627;
	#10 counter$count = 55628;
	#10 counter$count = 55629;
	#10 counter$count = 55630;
	#10 counter$count = 55631;
	#10 counter$count = 55632;
	#10 counter$count = 55633;
	#10 counter$count = 55634;
	#10 counter$count = 55635;
	#10 counter$count = 55636;
	#10 counter$count = 55637;
	#10 counter$count = 55638;
	#10 counter$count = 55639;
	#10 counter$count = 55640;
	#10 counter$count = 55641;
	#10 counter$count = 55642;
	#10 counter$count = 55643;
	#10 counter$count = 55644;
	#10 counter$count = 55645;
	#10 counter$count = 55646;
	#10 counter$count = 55647;
	#10 counter$count = 55648;
	#10 counter$count = 55649;
	#10 counter$count = 55650;
	#10 counter$count = 55651;
	#10 counter$count = 55652;
	#10 counter$count = 55653;
	#10 counter$count = 55654;
	#10 counter$count = 55655;
	#10 counter$count = 55656;
	#10 counter$count = 55657;
	#10 counter$count = 55658;
	#10 counter$count = 55659;
	#10 counter$count = 55660;
	#10 counter$count = 55661;
	#10 counter$count = 55662;
	#10 counter$count = 55663;
	#10 counter$count = 55664;
	#10 counter$count = 55665;
	#10 counter$count = 55666;
	#10 counter$count = 55667;
	#10 counter$count = 55668;
	#10 counter$count = 55669;
	#10 counter$count = 55670;
	#10 counter$count = 55671;
	#10 counter$count = 55672;
	#10 counter$count = 55673;
	#10 counter$count = 55674;
	#10 counter$count = 55675;
	#10 counter$count = 55676;
	#10 counter$count = 55677;
	#10 counter$count = 55678;
	#10 counter$count = 55679;
	#10 counter$count = 55680;
	#10 counter$count = 55681;
	#10 counter$count = 55682;
	#10 counter$count = 55683;
	#10 counter$count = 55684;
	#10 counter$count = 55685;
	#10 counter$count = 55686;
	#10 counter$count = 55687;
	#10 counter$count = 55688;
	#10 counter$count = 55689;
	#10 counter$count = 55690;
	#10 counter$count = 55691;
	#10 counter$count = 55692;
	#10 counter$count = 55693;
	#10 counter$count = 55694;
	#10 counter$count = 55695;
	#10 counter$count = 55696;
	#10 counter$count = 55697;
	#10 counter$count = 55698;
	#10 counter$count = 55699;
	#10 counter$count = 55700;
	#10 counter$count = 55701;
	#10 counter$count = 55702;
	#10 counter$count = 55703;
	#10 counter$count = 55704;
	#10 counter$count = 55705;
	#10 counter$count = 55706;
	#10 counter$count = 55707;
	#10 counter$count = 55708;
	#10 counter$count = 55709;
	#10 counter$count = 55710;
	#10 counter$count = 55711;
	#10 counter$count = 55712;
	#10 counter$count = 55713;
	#10 counter$count = 55714;
	#10 counter$count = 55715;
	#10 counter$count = 55716;
	#10 counter$count = 55717;
	#10 counter$count = 55718;
	#10 counter$count = 55719;
	#10 counter$count = 55720;
	#10 counter$count = 55721;
	#10 counter$count = 55722;
	#10 counter$count = 55723;
	#10 counter$count = 55724;
	#10 counter$count = 55725;
	#10 counter$count = 55726;
	#10 counter$count = 55727;
	#10 counter$count = 55728;
	#10 counter$count = 55729;
	#10 counter$count = 55730;
	#10 counter$count = 55731;
	#10 counter$count = 55732;
	#10 counter$count = 55733;
	#10 counter$count = 55734;
	#10 counter$count = 55735;
	#10 counter$count = 55736;
	#10 counter$count = 55737;
	#10 counter$count = 55738;
	#10 counter$count = 55739;
	#10 counter$count = 55740;
	#10 counter$count = 55741;
	#10 counter$count = 55742;
	#10 counter$count = 55743;
	#10 counter$count = 55744;
	#10 counter$count = 55745;
	#10 counter$count = 55746;
	#10 counter$count = 55747;
	#10 counter$count = 55748;
	#10 counter$count = 55749;
	#10 counter$count = 55750;
	#10 counter$count = 55751;
	#10 counter$count = 55752;
	#10 counter$count = 55753;
	#10 counter$count = 55754;
	#10 counter$count = 55755;
	#10 counter$count = 55756;
	#10 counter$count = 55757;
	#10 counter$count = 55758;
	#10 counter$count = 55759;
	#10 counter$count = 55760;
	#10 counter$count = 55761;
	#10 counter$count = 55762;
	#10 counter$count = 55763;
	#10 counter$count = 55764;
	#10 counter$count = 55765;
	#10 counter$count = 55766;
	#10 counter$count = 55767;
	#10 counter$count = 55768;
	#10 counter$count = 55769;
	#10 counter$count = 55770;
	#10 counter$count = 55771;
	#10 counter$count = 55772;
	#10 counter$count = 55773;
	#10 counter$count = 55774;
	#10 counter$count = 55775;
	#10 counter$count = 55776;
	#10 counter$count = 55777;
	#10 counter$count = 55778;
	#10 counter$count = 55779;
	#10 counter$count = 55780;
	#10 counter$count = 55781;
	#10 counter$count = 55782;
	#10 counter$count = 55783;
	#10 counter$count = 55784;
	#10 counter$count = 55785;
	#10 counter$count = 55786;
	#10 counter$count = 55787;
	#10 counter$count = 55788;
	#10 counter$count = 55789;
	#10 counter$count = 55790;
	#10 counter$count = 55791;
	#10 counter$count = 55792;
	#10 counter$count = 55793;
	#10 counter$count = 55794;
	#10 counter$count = 55795;
	#10 counter$count = 55796;
	#10 counter$count = 55797;
	#10 counter$count = 55798;
	#10 counter$count = 55799;
	#10 counter$count = 55800;
	#10 counter$count = 55801;
	#10 counter$count = 55802;
	#10 counter$count = 55803;
	#10 counter$count = 55804;
	#10 counter$count = 55805;
	#10 counter$count = 55806;
	#10 counter$count = 55807;
	#10 counter$count = 55808;
	#10 counter$count = 55809;
	#10 counter$count = 55810;
	#10 counter$count = 55811;
	#10 counter$count = 55812;
	#10 counter$count = 55813;
	#10 counter$count = 55814;
	#10 counter$count = 55815;
	#10 counter$count = 55816;
	#10 counter$count = 55817;
	#10 counter$count = 55818;
	#10 counter$count = 55819;
	#10 counter$count = 55820;
	#10 counter$count = 55821;
	#10 counter$count = 55822;
	#10 counter$count = 55823;
	#10 counter$count = 55824;
	#10 counter$count = 55825;
	#10 counter$count = 55826;
	#10 counter$count = 55827;
	#10 counter$count = 55828;
	#10 counter$count = 55829;
	#10 counter$count = 55830;
	#10 counter$count = 55831;
	#10 counter$count = 55832;
	#10 counter$count = 55833;
	#10 counter$count = 55834;
	#10 counter$count = 55835;
	#10 counter$count = 55836;
	#10 counter$count = 55837;
	#10 counter$count = 55838;
	#10 counter$count = 55839;
	#10 counter$count = 55840;
	#10 counter$count = 55841;
	#10 counter$count = 55842;
	#10 counter$count = 55843;
	#10 counter$count = 55844;
	#10 counter$count = 55845;
	#10 counter$count = 55846;
	#10 counter$count = 55847;
	#10 counter$count = 55848;
	#10 counter$count = 55849;
	#10 counter$count = 55850;
	#10 counter$count = 55851;
	#10 counter$count = 55852;
	#10 counter$count = 55853;
	#10 counter$count = 55854;
	#10 counter$count = 55855;
	#10 counter$count = 55856;
	#10 counter$count = 55857;
	#10 counter$count = 55858;
	#10 counter$count = 55859;
	#10 counter$count = 55860;
	#10 counter$count = 55861;
	#10 counter$count = 55862;
	#10 counter$count = 55863;
	#10 counter$count = 55864;
	#10 counter$count = 55865;
	#10 counter$count = 55866;
	#10 counter$count = 55867;
	#10 counter$count = 55868;
	#10 counter$count = 55869;
	#10 counter$count = 55870;
	#10 counter$count = 55871;
	#10 counter$count = 55872;
	#10 counter$count = 55873;
	#10 counter$count = 55874;
	#10 counter$count = 55875;
	#10 counter$count = 55876;
	#10 counter$count = 55877;
	#10 counter$count = 55878;
	#10 counter$count = 55879;
	#10 counter$count = 55880;
	#10 counter$count = 55881;
	#10 counter$count = 55882;
	#10 counter$count = 55883;
	#10 counter$count = 55884;
	#10 counter$count = 55885;
	#10 counter$count = 55886;
	#10 counter$count = 55887;
	#10 counter$count = 55888;
	#10 counter$count = 55889;
	#10 counter$count = 55890;
	#10 counter$count = 55891;
	#10 counter$count = 55892;
	#10 counter$count = 55893;
	#10 counter$count = 55894;
	#10 counter$count = 55895;
	#10 counter$count = 55896;
	#10 counter$count = 55897;
	#10 counter$count = 55898;
	#10 counter$count = 55899;
	#10 counter$count = 55900;
	#10 counter$count = 55901;
	#10 counter$count = 55902;
	#10 counter$count = 55903;
	#10 counter$count = 55904;
	#10 counter$count = 55905;
	#10 counter$count = 55906;
	#10 counter$count = 55907;
	#10 counter$count = 55908;
	#10 counter$count = 55909;
	#10 counter$count = 55910;
	#10 counter$count = 55911;
	#10 counter$count = 55912;
	#10 counter$count = 55913;
	#10 counter$count = 55914;
	#10 counter$count = 55915;
	#10 counter$count = 55916;
	#10 counter$count = 55917;
	#10 counter$count = 55918;
	#10 counter$count = 55919;
	#10 counter$count = 55920;
	#10 counter$count = 55921;
	#10 counter$count = 55922;
	#10 counter$count = 55923;
	#10 counter$count = 55924;
	#10 counter$count = 55925;
	#10 counter$count = 55926;
	#10 counter$count = 55927;
	#10 counter$count = 55928;
	#10 counter$count = 55929;
	#10 counter$count = 55930;
	#10 counter$count = 55931;
	#10 counter$count = 55932;
	#10 counter$count = 55933;
	#10 counter$count = 55934;
	#10 counter$count = 55935;
	#10 counter$count = 55936;
	#10 counter$count = 55937;
	#10 counter$count = 55938;
	#10 counter$count = 55939;
	#10 counter$count = 55940;
	#10 counter$count = 55941;
	#10 counter$count = 55942;
	#10 counter$count = 55943;
	#10 counter$count = 55944;
	#10 counter$count = 55945;
	#10 counter$count = 55946;
	#10 counter$count = 55947;
	#10 counter$count = 55948;
	#10 counter$count = 55949;
	#10 counter$count = 55950;
	#10 counter$count = 55951;
	#10 counter$count = 55952;
	#10 counter$count = 55953;
	#10 counter$count = 55954;
	#10 counter$count = 55955;
	#10 counter$count = 55956;
	#10 counter$count = 55957;
	#10 counter$count = 55958;
	#10 counter$count = 55959;
	#10 counter$count = 55960;
	#10 counter$count = 55961;
	#10 counter$count = 55962;
	#10 counter$count = 55963;
	#10 counter$count = 55964;
	#10 counter$count = 55965;
	#10 counter$count = 55966;
	#10 counter$count = 55967;
	#10 counter$count = 55968;
	#10 counter$count = 55969;
	#10 counter$count = 55970;
	#10 counter$count = 55971;
	#10 counter$count = 55972;
	#10 counter$count = 55973;
	#10 counter$count = 55974;
	#10 counter$count = 55975;
	#10 counter$count = 55976;
	#10 counter$count = 55977;
	#10 counter$count = 55978;
	#10 counter$count = 55979;
	#10 counter$count = 55980;
	#10 counter$count = 55981;
	#10 counter$count = 55982;
	#10 counter$count = 55983;
	#10 counter$count = 55984;
	#10 counter$count = 55985;
	#10 counter$count = 55986;
	#10 counter$count = 55987;
	#10 counter$count = 55988;
	#10 counter$count = 55989;
	#10 counter$count = 55990;
	#10 counter$count = 55991;
	#10 counter$count = 55992;
	#10 counter$count = 55993;
	#10 counter$count = 55994;
	#10 counter$count = 55995;
	#10 counter$count = 55996;
	#10 counter$count = 55997;
	#10 counter$count = 55998;
	#10 counter$count = 55999;
	#10 counter$count = 56000;
	#10 counter$count = 56001;
	#10 counter$count = 56002;
	#10 counter$count = 56003;
	#10 counter$count = 56004;
	#10 counter$count = 56005;
	#10 counter$count = 56006;
	#10 counter$count = 56007;
	#10 counter$count = 56008;
	#10 counter$count = 56009;
	#10 counter$count = 56010;
	#10 counter$count = 56011;
	#10 counter$count = 56012;
	#10 counter$count = 56013;
	#10 counter$count = 56014;
	#10 counter$count = 56015;
	#10 counter$count = 56016;
	#10 counter$count = 56017;
	#10 counter$count = 56018;
	#10 counter$count = 56019;
	#10 counter$count = 56020;
	#10 counter$count = 56021;
	#10 counter$count = 56022;
	#10 counter$count = 56023;
	#10 counter$count = 56024;
	#10 counter$count = 56025;
	#10 counter$count = 56026;
	#10 counter$count = 56027;
	#10 counter$count = 56028;
	#10 counter$count = 56029;
	#10 counter$count = 56030;
	#10 counter$count = 56031;
	#10 counter$count = 56032;
	#10 counter$count = 56033;
	#10 counter$count = 56034;
	#10 counter$count = 56035;
	#10 counter$count = 56036;
	#10 counter$count = 56037;
	#10 counter$count = 56038;
	#10 counter$count = 56039;
	#10 counter$count = 56040;
	#10 counter$count = 56041;
	#10 counter$count = 56042;
	#10 counter$count = 56043;
	#10 counter$count = 56044;
	#10 counter$count = 56045;
	#10 counter$count = 56046;
	#10 counter$count = 56047;
	#10 counter$count = 56048;
	#10 counter$count = 56049;
	#10 counter$count = 56050;
	#10 counter$count = 56051;
	#10 counter$count = 56052;
	#10 counter$count = 56053;
	#10 counter$count = 56054;
	#10 counter$count = 56055;
	#10 counter$count = 56056;
	#10 counter$count = 56057;
	#10 counter$count = 56058;
	#10 counter$count = 56059;
	#10 counter$count = 56060;
	#10 counter$count = 56061;
	#10 counter$count = 56062;
	#10 counter$count = 56063;
	#10 counter$count = 56064;
	#10 counter$count = 56065;
	#10 counter$count = 56066;
	#10 counter$count = 56067;
	#10 counter$count = 56068;
	#10 counter$count = 56069;
	#10 counter$count = 56070;
	#10 counter$count = 56071;
	#10 counter$count = 56072;
	#10 counter$count = 56073;
	#10 counter$count = 56074;
	#10 counter$count = 56075;
	#10 counter$count = 56076;
	#10 counter$count = 56077;
	#10 counter$count = 56078;
	#10 counter$count = 56079;
	#10 counter$count = 56080;
	#10 counter$count = 56081;
	#10 counter$count = 56082;
	#10 counter$count = 56083;
	#10 counter$count = 56084;
	#10 counter$count = 56085;
	#10 counter$count = 56086;
	#10 counter$count = 56087;
	#10 counter$count = 56088;
	#10 counter$count = 56089;
	#10 counter$count = 56090;
	#10 counter$count = 56091;
	#10 counter$count = 56092;
	#10 counter$count = 56093;
	#10 counter$count = 56094;
	#10 counter$count = 56095;
	#10 counter$count = 56096;
	#10 counter$count = 56097;
	#10 counter$count = 56098;
	#10 counter$count = 56099;
	#10 counter$count = 56100;
	#10 counter$count = 56101;
	#10 counter$count = 56102;
	#10 counter$count = 56103;
	#10 counter$count = 56104;
	#10 counter$count = 56105;
	#10 counter$count = 56106;
	#10 counter$count = 56107;
	#10 counter$count = 56108;
	#10 counter$count = 56109;
	#10 counter$count = 56110;
	#10 counter$count = 56111;
	#10 counter$count = 56112;
	#10 counter$count = 56113;
	#10 counter$count = 56114;
	#10 counter$count = 56115;
	#10 counter$count = 56116;
	#10 counter$count = 56117;
	#10 counter$count = 56118;
	#10 counter$count = 56119;
	#10 counter$count = 56120;
	#10 counter$count = 56121;
	#10 counter$count = 56122;
	#10 counter$count = 56123;
	#10 counter$count = 56124;
	#10 counter$count = 56125;
	#10 counter$count = 56126;
	#10 counter$count = 56127;
	#10 counter$count = 56128;
	#10 counter$count = 56129;
	#10 counter$count = 56130;
	#10 counter$count = 56131;
	#10 counter$count = 56132;
	#10 counter$count = 56133;
	#10 counter$count = 56134;
	#10 counter$count = 56135;
	#10 counter$count = 56136;
	#10 counter$count = 56137;
	#10 counter$count = 56138;
	#10 counter$count = 56139;
	#10 counter$count = 56140;
	#10 counter$count = 56141;
	#10 counter$count = 56142;
	#10 counter$count = 56143;
	#10 counter$count = 56144;
	#10 counter$count = 56145;
	#10 counter$count = 56146;
	#10 counter$count = 56147;
	#10 counter$count = 56148;
	#10 counter$count = 56149;
	#10 counter$count = 56150;
	#10 counter$count = 56151;
	#10 counter$count = 56152;
	#10 counter$count = 56153;
	#10 counter$count = 56154;
	#10 counter$count = 56155;
	#10 counter$count = 56156;
	#10 counter$count = 56157;
	#10 counter$count = 56158;
	#10 counter$count = 56159;
	#10 counter$count = 56160;
	#10 counter$count = 56161;
	#10 counter$count = 56162;
	#10 counter$count = 56163;
	#10 counter$count = 56164;
	#10 counter$count = 56165;
	#10 counter$count = 56166;
	#10 counter$count = 56167;
	#10 counter$count = 56168;
	#10 counter$count = 56169;
	#10 counter$count = 56170;
	#10 counter$count = 56171;
	#10 counter$count = 56172;
	#10 counter$count = 56173;
	#10 counter$count = 56174;
	#10 counter$count = 56175;
	#10 counter$count = 56176;
	#10 counter$count = 56177;
	#10 counter$count = 56178;
	#10 counter$count = 56179;
	#10 counter$count = 56180;
	#10 counter$count = 56181;
	#10 counter$count = 56182;
	#10 counter$count = 56183;
	#10 counter$count = 56184;
	#10 counter$count = 56185;
	#10 counter$count = 56186;
	#10 counter$count = 56187;
	#10 counter$count = 56188;
	#10 counter$count = 56189;
	#10 counter$count = 56190;
	#10 counter$count = 56191;
	#10 counter$count = 56192;
	#10 counter$count = 56193;
	#10 counter$count = 56194;
	#10 counter$count = 56195;
	#10 counter$count = 56196;
	#10 counter$count = 56197;
	#10 counter$count = 56198;
	#10 counter$count = 56199;
	#10 counter$count = 56200;
	#10 counter$count = 56201;
	#10 counter$count = 56202;
	#10 counter$count = 56203;
	#10 counter$count = 56204;
	#10 counter$count = 56205;
	#10 counter$count = 56206;
	#10 counter$count = 56207;
	#10 counter$count = 56208;
	#10 counter$count = 56209;
	#10 counter$count = 56210;
	#10 counter$count = 56211;
	#10 counter$count = 56212;
	#10 counter$count = 56213;
	#10 counter$count = 56214;
	#10 counter$count = 56215;
	#10 counter$count = 56216;
	#10 counter$count = 56217;
	#10 counter$count = 56218;
	#10 counter$count = 56219;
	#10 counter$count = 56220;
	#10 counter$count = 56221;
	#10 counter$count = 56222;
	#10 counter$count = 56223;
	#10 counter$count = 56224;
	#10 counter$count = 56225;
	#10 counter$count = 56226;
	#10 counter$count = 56227;
	#10 counter$count = 56228;
	#10 counter$count = 56229;
	#10 counter$count = 56230;
	#10 counter$count = 56231;
	#10 counter$count = 56232;
	#10 counter$count = 56233;
	#10 counter$count = 56234;
	#10 counter$count = 56235;
	#10 counter$count = 56236;
	#10 counter$count = 56237;
	#10 counter$count = 56238;
	#10 counter$count = 56239;
	#10 counter$count = 56240;
	#10 counter$count = 56241;
	#10 counter$count = 56242;
	#10 counter$count = 56243;
	#10 counter$count = 56244;
	#10 counter$count = 56245;
	#10 counter$count = 56246;
	#10 counter$count = 56247;
	#10 counter$count = 56248;
	#10 counter$count = 56249;
	#10 counter$count = 56250;
	#10 counter$count = 56251;
	#10 counter$count = 56252;
	#10 counter$count = 56253;
	#10 counter$count = 56254;
	#10 counter$count = 56255;
	#10 counter$count = 56256;
	#10 counter$count = 56257;
	#10 counter$count = 56258;
	#10 counter$count = 56259;
	#10 counter$count = 56260;
	#10 counter$count = 56261;
	#10 counter$count = 56262;
	#10 counter$count = 56263;
	#10 counter$count = 56264;
	#10 counter$count = 56265;
	#10 counter$count = 56266;
	#10 counter$count = 56267;
	#10 counter$count = 56268;
	#10 counter$count = 56269;
	#10 counter$count = 56270;
	#10 counter$count = 56271;
	#10 counter$count = 56272;
	#10 counter$count = 56273;
	#10 counter$count = 56274;
	#10 counter$count = 56275;
	#10 counter$count = 56276;
	#10 counter$count = 56277;
	#10 counter$count = 56278;
	#10 counter$count = 56279;
	#10 counter$count = 56280;
	#10 counter$count = 56281;
	#10 counter$count = 56282;
	#10 counter$count = 56283;
	#10 counter$count = 56284;
	#10 counter$count = 56285;
	#10 counter$count = 56286;
	#10 counter$count = 56287;
	#10 counter$count = 56288;
	#10 counter$count = 56289;
	#10 counter$count = 56290;
	#10 counter$count = 56291;
	#10 counter$count = 56292;
	#10 counter$count = 56293;
	#10 counter$count = 56294;
	#10 counter$count = 56295;
	#10 counter$count = 56296;
	#10 counter$count = 56297;
	#10 counter$count = 56298;
	#10 counter$count = 56299;
	#10 counter$count = 56300;
	#10 counter$count = 56301;
	#10 counter$count = 56302;
	#10 counter$count = 56303;
	#10 counter$count = 56304;
	#10 counter$count = 56305;
	#10 counter$count = 56306;
	#10 counter$count = 56307;
	#10 counter$count = 56308;
	#10 counter$count = 56309;
	#10 counter$count = 56310;
	#10 counter$count = 56311;
	#10 counter$count = 56312;
	#10 counter$count = 56313;
	#10 counter$count = 56314;
	#10 counter$count = 56315;
	#10 counter$count = 56316;
	#10 counter$count = 56317;
	#10 counter$count = 56318;
	#10 counter$count = 56319;
	#10 counter$count = 56320;
	#10 counter$count = 56321;
	#10 counter$count = 56322;
	#10 counter$count = 56323;
	#10 counter$count = 56324;
	#10 counter$count = 56325;
	#10 counter$count = 56326;
	#10 counter$count = 56327;
	#10 counter$count = 56328;
	#10 counter$count = 56329;
	#10 counter$count = 56330;
	#10 counter$count = 56331;
	#10 counter$count = 56332;
	#10 counter$count = 56333;
	#10 counter$count = 56334;
	#10 counter$count = 56335;
	#10 counter$count = 56336;
	#10 counter$count = 56337;
	#10 counter$count = 56338;
	#10 counter$count = 56339;
	#10 counter$count = 56340;
	#10 counter$count = 56341;
	#10 counter$count = 56342;
	#10 counter$count = 56343;
	#10 counter$count = 56344;
	#10 counter$count = 56345;
	#10 counter$count = 56346;
	#10 counter$count = 56347;
	#10 counter$count = 56348;
	#10 counter$count = 56349;
	#10 counter$count = 56350;
	#10 counter$count = 56351;
	#10 counter$count = 56352;
	#10 counter$count = 56353;
	#10 counter$count = 56354;
	#10 counter$count = 56355;
	#10 counter$count = 56356;
	#10 counter$count = 56357;
	#10 counter$count = 56358;
	#10 counter$count = 56359;
	#10 counter$count = 56360;
	#10 counter$count = 56361;
	#10 counter$count = 56362;
	#10 counter$count = 56363;
	#10 counter$count = 56364;
	#10 counter$count = 56365;
	#10 counter$count = 56366;
	#10 counter$count = 56367;
	#10 counter$count = 56368;
	#10 counter$count = 56369;
	#10 counter$count = 56370;
	#10 counter$count = 56371;
	#10 counter$count = 56372;
	#10 counter$count = 56373;
	#10 counter$count = 56374;
	#10 counter$count = 56375;
	#10 counter$count = 56376;
	#10 counter$count = 56377;
	#10 counter$count = 56378;
	#10 counter$count = 56379;
	#10 counter$count = 56380;
	#10 counter$count = 56381;
	#10 counter$count = 56382;
	#10 counter$count = 56383;
	#10 counter$count = 56384;
	#10 counter$count = 56385;
	#10 counter$count = 56386;
	#10 counter$count = 56387;
	#10 counter$count = 56388;
	#10 counter$count = 56389;
	#10 counter$count = 56390;
	#10 counter$count = 56391;
	#10 counter$count = 56392;
	#10 counter$count = 56393;
	#10 counter$count = 56394;
	#10 counter$count = 56395;
	#10 counter$count = 56396;
	#10 counter$count = 56397;
	#10 counter$count = 56398;
	#10 counter$count = 56399;
	#10 counter$count = 56400;
	#10 counter$count = 56401;
	#10 counter$count = 56402;
	#10 counter$count = 56403;
	#10 counter$count = 56404;
	#10 counter$count = 56405;
	#10 counter$count = 56406;
	#10 counter$count = 56407;
	#10 counter$count = 56408;
	#10 counter$count = 56409;
	#10 counter$count = 56410;
	#10 counter$count = 56411;
	#10 counter$count = 56412;
	#10 counter$count = 56413;
	#10 counter$count = 56414;
	#10 counter$count = 56415;
	#10 counter$count = 56416;
	#10 counter$count = 56417;
	#10 counter$count = 56418;
	#10 counter$count = 56419;
	#10 counter$count = 56420;
	#10 counter$count = 56421;
	#10 counter$count = 56422;
	#10 counter$count = 56423;
	#10 counter$count = 56424;
	#10 counter$count = 56425;
	#10 counter$count = 56426;
	#10 counter$count = 56427;
	#10 counter$count = 56428;
	#10 counter$count = 56429;
	#10 counter$count = 56430;
	#10 counter$count = 56431;
	#10 counter$count = 56432;
	#10 counter$count = 56433;
	#10 counter$count = 56434;
	#10 counter$count = 56435;
	#10 counter$count = 56436;
	#10 counter$count = 56437;
	#10 counter$count = 56438;
	#10 counter$count = 56439;
	#10 counter$count = 56440;
	#10 counter$count = 56441;
	#10 counter$count = 56442;
	#10 counter$count = 56443;
	#10 counter$count = 56444;
	#10 counter$count = 56445;
	#10 counter$count = 56446;
	#10 counter$count = 56447;
	#10 counter$count = 56448;
	#10 counter$count = 56449;
	#10 counter$count = 56450;
	#10 counter$count = 56451;
	#10 counter$count = 56452;
	#10 counter$count = 56453;
	#10 counter$count = 56454;
	#10 counter$count = 56455;
	#10 counter$count = 56456;
	#10 counter$count = 56457;
	#10 counter$count = 56458;
	#10 counter$count = 56459;
	#10 counter$count = 56460;
	#10 counter$count = 56461;
	#10 counter$count = 56462;
	#10 counter$count = 56463;
	#10 counter$count = 56464;
	#10 counter$count = 56465;
	#10 counter$count = 56466;
	#10 counter$count = 56467;
	#10 counter$count = 56468;
	#10 counter$count = 56469;
	#10 counter$count = 56470;
	#10 counter$count = 56471;
	#10 counter$count = 56472;
	#10 counter$count = 56473;
	#10 counter$count = 56474;
	#10 counter$count = 56475;
	#10 counter$count = 56476;
	#10 counter$count = 56477;
	#10 counter$count = 56478;
	#10 counter$count = 56479;
	#10 counter$count = 56480;
	#10 counter$count = 56481;
	#10 counter$count = 56482;
	#10 counter$count = 56483;
	#10 counter$count = 56484;
	#10 counter$count = 56485;
	#10 counter$count = 56486;
	#10 counter$count = 56487;
	#10 counter$count = 56488;
	#10 counter$count = 56489;
	#10 counter$count = 56490;
	#10 counter$count = 56491;
	#10 counter$count = 56492;
	#10 counter$count = 56493;
	#10 counter$count = 56494;
	#10 counter$count = 56495;
	#10 counter$count = 56496;
	#10 counter$count = 56497;
	#10 counter$count = 56498;
	#10 counter$count = 56499;
	#10 counter$count = 56500;
	#10 counter$count = 56501;
	#10 counter$count = 56502;
	#10 counter$count = 56503;
	#10 counter$count = 56504;
	#10 counter$count = 56505;
	#10 counter$count = 56506;
	#10 counter$count = 56507;
	#10 counter$count = 56508;
	#10 counter$count = 56509;
	#10 counter$count = 56510;
	#10 counter$count = 56511;
	#10 counter$count = 56512;
	#10 counter$count = 56513;
	#10 counter$count = 56514;
	#10 counter$count = 56515;
	#10 counter$count = 56516;
	#10 counter$count = 56517;
	#10 counter$count = 56518;
	#10 counter$count = 56519;
	#10 counter$count = 56520;
	#10 counter$count = 56521;
	#10 counter$count = 56522;
	#10 counter$count = 56523;
	#10 counter$count = 56524;
	#10 counter$count = 56525;
	#10 counter$count = 56526;
	#10 counter$count = 56527;
	#10 counter$count = 56528;
	#10 counter$count = 56529;
	#10 counter$count = 56530;
	#10 counter$count = 56531;
	#10 counter$count = 56532;
	#10 counter$count = 56533;
	#10 counter$count = 56534;
	#10 counter$count = 56535;
	#10 counter$count = 56536;
	#10 counter$count = 56537;
	#10 counter$count = 56538;
	#10 counter$count = 56539;
	#10 counter$count = 56540;
	#10 counter$count = 56541;
	#10 counter$count = 56542;
	#10 counter$count = 56543;
	#10 counter$count = 56544;
	#10 counter$count = 56545;
	#10 counter$count = 56546;
	#10 counter$count = 56547;
	#10 counter$count = 56548;
	#10 counter$count = 56549;
	#10 counter$count = 56550;
	#10 counter$count = 56551;
	#10 counter$count = 56552;
	#10 counter$count = 56553;
	#10 counter$count = 56554;
	#10 counter$count = 56555;
	#10 counter$count = 56556;
	#10 counter$count = 56557;
	#10 counter$count = 56558;
	#10 counter$count = 56559;
	#10 counter$count = 56560;
	#10 counter$count = 56561;
	#10 counter$count = 56562;
	#10 counter$count = 56563;
	#10 counter$count = 56564;
	#10 counter$count = 56565;
	#10 counter$count = 56566;
	#10 counter$count = 56567;
	#10 counter$count = 56568;
	#10 counter$count = 56569;
	#10 counter$count = 56570;
	#10 counter$count = 56571;
	#10 counter$count = 56572;
	#10 counter$count = 56573;
	#10 counter$count = 56574;
	#10 counter$count = 56575;
	#10 counter$count = 56576;
	#10 counter$count = 56577;
	#10 counter$count = 56578;
	#10 counter$count = 56579;
	#10 counter$count = 56580;
	#10 counter$count = 56581;
	#10 counter$count = 56582;
	#10 counter$count = 56583;
	#10 counter$count = 56584;
	#10 counter$count = 56585;
	#10 counter$count = 56586;
	#10 counter$count = 56587;
	#10 counter$count = 56588;
	#10 counter$count = 56589;
	#10 counter$count = 56590;
	#10 counter$count = 56591;
	#10 counter$count = 56592;
	#10 counter$count = 56593;
	#10 counter$count = 56594;
	#10 counter$count = 56595;
	#10 counter$count = 56596;
	#10 counter$count = 56597;
	#10 counter$count = 56598;
	#10 counter$count = 56599;
	#10 counter$count = 56600;
	#10 counter$count = 56601;
	#10 counter$count = 56602;
	#10 counter$count = 56603;
	#10 counter$count = 56604;
	#10 counter$count = 56605;
	#10 counter$count = 56606;
	#10 counter$count = 56607;
	#10 counter$count = 56608;
	#10 counter$count = 56609;
	#10 counter$count = 56610;
	#10 counter$count = 56611;
	#10 counter$count = 56612;
	#10 counter$count = 56613;
	#10 counter$count = 56614;
	#10 counter$count = 56615;
	#10 counter$count = 56616;
	#10 counter$count = 56617;
	#10 counter$count = 56618;
	#10 counter$count = 56619;
	#10 counter$count = 56620;
	#10 counter$count = 56621;
	#10 counter$count = 56622;
	#10 counter$count = 56623;
	#10 counter$count = 56624;
	#10 counter$count = 56625;
	#10 counter$count = 56626;
	#10 counter$count = 56627;
	#10 counter$count = 56628;
	#10 counter$count = 56629;
	#10 counter$count = 56630;
	#10 counter$count = 56631;
	#10 counter$count = 56632;
	#10 counter$count = 56633;
	#10 counter$count = 56634;
	#10 counter$count = 56635;
	#10 counter$count = 56636;
	#10 counter$count = 56637;
	#10 counter$count = 56638;
	#10 counter$count = 56639;
	#10 counter$count = 56640;
	#10 counter$count = 56641;
	#10 counter$count = 56642;
	#10 counter$count = 56643;
	#10 counter$count = 56644;
	#10 counter$count = 56645;
	#10 counter$count = 56646;
	#10 counter$count = 56647;
	#10 counter$count = 56648;
	#10 counter$count = 56649;
	#10 counter$count = 56650;
	#10 counter$count = 56651;
	#10 counter$count = 56652;
	#10 counter$count = 56653;
	#10 counter$count = 56654;
	#10 counter$count = 56655;
	#10 counter$count = 56656;
	#10 counter$count = 56657;
	#10 counter$count = 56658;
	#10 counter$count = 56659;
	#10 counter$count = 56660;
	#10 counter$count = 56661;
	#10 counter$count = 56662;
	#10 counter$count = 56663;
	#10 counter$count = 56664;
	#10 counter$count = 56665;
	#10 counter$count = 56666;
	#10 counter$count = 56667;
	#10 counter$count = 56668;
	#10 counter$count = 56669;
	#10 counter$count = 56670;
	#10 counter$count = 56671;
	#10 counter$count = 56672;
	#10 counter$count = 56673;
	#10 counter$count = 56674;
	#10 counter$count = 56675;
	#10 counter$count = 56676;
	#10 counter$count = 56677;
	#10 counter$count = 56678;
	#10 counter$count = 56679;
	#10 counter$count = 56680;
	#10 counter$count = 56681;
	#10 counter$count = 56682;
	#10 counter$count = 56683;
	#10 counter$count = 56684;
	#10 counter$count = 56685;
	#10 counter$count = 56686;
	#10 counter$count = 56687;
	#10 counter$count = 56688;
	#10 counter$count = 56689;
	#10 counter$count = 56690;
	#10 counter$count = 56691;
	#10 counter$count = 56692;
	#10 counter$count = 56693;
	#10 counter$count = 56694;
	#10 counter$count = 56695;
	#10 counter$count = 56696;
	#10 counter$count = 56697;
	#10 counter$count = 56698;
	#10 counter$count = 56699;
	#10 counter$count = 56700;
	#10 counter$count = 56701;
	#10 counter$count = 56702;
	#10 counter$count = 56703;
	#10 counter$count = 56704;
	#10 counter$count = 56705;
	#10 counter$count = 56706;
	#10 counter$count = 56707;
	#10 counter$count = 56708;
	#10 counter$count = 56709;
	#10 counter$count = 56710;
	#10 counter$count = 56711;
	#10 counter$count = 56712;
	#10 counter$count = 56713;
	#10 counter$count = 56714;
	#10 counter$count = 56715;
	#10 counter$count = 56716;
	#10 counter$count = 56717;
	#10 counter$count = 56718;
	#10 counter$count = 56719;
	#10 counter$count = 56720;
	#10 counter$count = 56721;
	#10 counter$count = 56722;
	#10 counter$count = 56723;
	#10 counter$count = 56724;
	#10 counter$count = 56725;
	#10 counter$count = 56726;
	#10 counter$count = 56727;
	#10 counter$count = 56728;
	#10 counter$count = 56729;
	#10 counter$count = 56730;
	#10 counter$count = 56731;
	#10 counter$count = 56732;
	#10 counter$count = 56733;
	#10 counter$count = 56734;
	#10 counter$count = 56735;
	#10 counter$count = 56736;
	#10 counter$count = 56737;
	#10 counter$count = 56738;
	#10 counter$count = 56739;
	#10 counter$count = 56740;
	#10 counter$count = 56741;
	#10 counter$count = 56742;
	#10 counter$count = 56743;
	#10 counter$count = 56744;
	#10 counter$count = 56745;
	#10 counter$count = 56746;
	#10 counter$count = 56747;
	#10 counter$count = 56748;
	#10 counter$count = 56749;
	#10 counter$count = 56750;
	#10 counter$count = 56751;
	#10 counter$count = 56752;
	#10 counter$count = 56753;
	#10 counter$count = 56754;
	#10 counter$count = 56755;
	#10 counter$count = 56756;
	#10 counter$count = 56757;
	#10 counter$count = 56758;
	#10 counter$count = 56759;
	#10 counter$count = 56760;
	#10 counter$count = 56761;
	#10 counter$count = 56762;
	#10 counter$count = 56763;
	#10 counter$count = 56764;
	#10 counter$count = 56765;
	#10 counter$count = 56766;
	#10 counter$count = 56767;
	#10 counter$count = 56768;
	#10 counter$count = 56769;
	#10 counter$count = 56770;
	#10 counter$count = 56771;
	#10 counter$count = 56772;
	#10 counter$count = 56773;
	#10 counter$count = 56774;
	#10 counter$count = 56775;
	#10 counter$count = 56776;
	#10 counter$count = 56777;
	#10 counter$count = 56778;
	#10 counter$count = 56779;
	#10 counter$count = 56780;
	#10 counter$count = 56781;
	#10 counter$count = 56782;
	#10 counter$count = 56783;
	#10 counter$count = 56784;
	#10 counter$count = 56785;
	#10 counter$count = 56786;
	#10 counter$count = 56787;
	#10 counter$count = 56788;
	#10 counter$count = 56789;
	#10 counter$count = 56790;
	#10 counter$count = 56791;
	#10 counter$count = 56792;
	#10 counter$count = 56793;
	#10 counter$count = 56794;
	#10 counter$count = 56795;
	#10 counter$count = 56796;
	#10 counter$count = 56797;
	#10 counter$count = 56798;
	#10 counter$count = 56799;
	#10 counter$count = 56800;
	#10 counter$count = 56801;
	#10 counter$count = 56802;
	#10 counter$count = 56803;
	#10 counter$count = 56804;
	#10 counter$count = 56805;
	#10 counter$count = 56806;
	#10 counter$count = 56807;
	#10 counter$count = 56808;
	#10 counter$count = 56809;
	#10 counter$count = 56810;
	#10 counter$count = 56811;
	#10 counter$count = 56812;
	#10 counter$count = 56813;
	#10 counter$count = 56814;
	#10 counter$count = 56815;
	#10 counter$count = 56816;
	#10 counter$count = 56817;
	#10 counter$count = 56818;
	#10 counter$count = 56819;
	#10 counter$count = 56820;
	#10 counter$count = 56821;
	#10 counter$count = 56822;
	#10 counter$count = 56823;
	#10 counter$count = 56824;
	#10 counter$count = 56825;
	#10 counter$count = 56826;
	#10 counter$count = 56827;
	#10 counter$count = 56828;
	#10 counter$count = 56829;
	#10 counter$count = 56830;
	#10 counter$count = 56831;
	#10 counter$count = 56832;
	#10 counter$count = 56833;
	#10 counter$count = 56834;
	#10 counter$count = 56835;
	#10 counter$count = 56836;
	#10 counter$count = 56837;
	#10 counter$count = 56838;
	#10 counter$count = 56839;
	#10 counter$count = 56840;
	#10 counter$count = 56841;
	#10 counter$count = 56842;
	#10 counter$count = 56843;
	#10 counter$count = 56844;
	#10 counter$count = 56845;
	#10 counter$count = 56846;
	#10 counter$count = 56847;
	#10 counter$count = 56848;
	#10 counter$count = 56849;
	#10 counter$count = 56850;
	#10 counter$count = 56851;
	#10 counter$count = 56852;
	#10 counter$count = 56853;
	#10 counter$count = 56854;
	#10 counter$count = 56855;
	#10 counter$count = 56856;
	#10 counter$count = 56857;
	#10 counter$count = 56858;
	#10 counter$count = 56859;
	#10 counter$count = 56860;
	#10 counter$count = 56861;
	#10 counter$count = 56862;
	#10 counter$count = 56863;
	#10 counter$count = 56864;
	#10 counter$count = 56865;
	#10 counter$count = 56866;
	#10 counter$count = 56867;
	#10 counter$count = 56868;
	#10 counter$count = 56869;
	#10 counter$count = 56870;
	#10 counter$count = 56871;
	#10 counter$count = 56872;
	#10 counter$count = 56873;
	#10 counter$count = 56874;
	#10 counter$count = 56875;
	#10 counter$count = 56876;
	#10 counter$count = 56877;
	#10 counter$count = 56878;
	#10 counter$count = 56879;
	#10 counter$count = 56880;
	#10 counter$count = 56881;
	#10 counter$count = 56882;
	#10 counter$count = 56883;
	#10 counter$count = 56884;
	#10 counter$count = 56885;
	#10 counter$count = 56886;
	#10 counter$count = 56887;
	#10 counter$count = 56888;
	#10 counter$count = 56889;
	#10 counter$count = 56890;
	#10 counter$count = 56891;
	#10 counter$count = 56892;
	#10 counter$count = 56893;
	#10 counter$count = 56894;
	#10 counter$count = 56895;
	#10 counter$count = 56896;
	#10 counter$count = 56897;
	#10 counter$count = 56898;
	#10 counter$count = 56899;
	#10 counter$count = 56900;
	#10 counter$count = 56901;
	#10 counter$count = 56902;
	#10 counter$count = 56903;
	#10 counter$count = 56904;
	#10 counter$count = 56905;
	#10 counter$count = 56906;
	#10 counter$count = 56907;
	#10 counter$count = 56908;
	#10 counter$count = 56909;
	#10 counter$count = 56910;
	#10 counter$count = 56911;
	#10 counter$count = 56912;
	#10 counter$count = 56913;
	#10 counter$count = 56914;
	#10 counter$count = 56915;
	#10 counter$count = 56916;
	#10 counter$count = 56917;
	#10 counter$count = 56918;
	#10 counter$count = 56919;
	#10 counter$count = 56920;
	#10 counter$count = 56921;
	#10 counter$count = 56922;
	#10 counter$count = 56923;
	#10 counter$count = 56924;
	#10 counter$count = 56925;
	#10 counter$count = 56926;
	#10 counter$count = 56927;
	#10 counter$count = 56928;
	#10 counter$count = 56929;
	#10 counter$count = 56930;
	#10 counter$count = 56931;
	#10 counter$count = 56932;
	#10 counter$count = 56933;
	#10 counter$count = 56934;
	#10 counter$count = 56935;
	#10 counter$count = 56936;
	#10 counter$count = 56937;
	#10 counter$count = 56938;
	#10 counter$count = 56939;
	#10 counter$count = 56940;
	#10 counter$count = 56941;
	#10 counter$count = 56942;
	#10 counter$count = 56943;
	#10 counter$count = 56944;
	#10 counter$count = 56945;
	#10 counter$count = 56946;
	#10 counter$count = 56947;
	#10 counter$count = 56948;
	#10 counter$count = 56949;
	#10 counter$count = 56950;
	#10 counter$count = 56951;
	#10 counter$count = 56952;
	#10 counter$count = 56953;
	#10 counter$count = 56954;
	#10 counter$count = 56955;
	#10 counter$count = 56956;
	#10 counter$count = 56957;
	#10 counter$count = 56958;
	#10 counter$count = 56959;
	#10 counter$count = 56960;
	#10 counter$count = 56961;
	#10 counter$count = 56962;
	#10 counter$count = 56963;
	#10 counter$count = 56964;
	#10 counter$count = 56965;
	#10 counter$count = 56966;
	#10 counter$count = 56967;
	#10 counter$count = 56968;
	#10 counter$count = 56969;
	#10 counter$count = 56970;
	#10 counter$count = 56971;
	#10 counter$count = 56972;
	#10 counter$count = 56973;
	#10 counter$count = 56974;
	#10 counter$count = 56975;
	#10 counter$count = 56976;
	#10 counter$count = 56977;
	#10 counter$count = 56978;
	#10 counter$count = 56979;
	#10 counter$count = 56980;
	#10 counter$count = 56981;
	#10 counter$count = 56982;
	#10 counter$count = 56983;
	#10 counter$count = 56984;
	#10 counter$count = 56985;
	#10 counter$count = 56986;
	#10 counter$count = 56987;
	#10 counter$count = 56988;
	#10 counter$count = 56989;
	#10 counter$count = 56990;
	#10 counter$count = 56991;
	#10 counter$count = 56992;
	#10 counter$count = 56993;
	#10 counter$count = 56994;
	#10 counter$count = 56995;
	#10 counter$count = 56996;
	#10 counter$count = 56997;
	#10 counter$count = 56998;
	#10 counter$count = 56999;
	#10 counter$count = 57000;
	#10 counter$count = 57001;
	#10 counter$count = 57002;
	#10 counter$count = 57003;
	#10 counter$count = 57004;
	#10 counter$count = 57005;
	#10 counter$count = 57006;
	#10 counter$count = 57007;
	#10 counter$count = 57008;
	#10 counter$count = 57009;
	#10 counter$count = 57010;
	#10 counter$count = 57011;
	#10 counter$count = 57012;
	#10 counter$count = 57013;
	#10 counter$count = 57014;
	#10 counter$count = 57015;
	#10 counter$count = 57016;
	#10 counter$count = 57017;
	#10 counter$count = 57018;
	#10 counter$count = 57019;
	#10 counter$count = 57020;
	#10 counter$count = 57021;
	#10 counter$count = 57022;
	#10 counter$count = 57023;
	#10 counter$count = 57024;
	#10 counter$count = 57025;
	#10 counter$count = 57026;
	#10 counter$count = 57027;
	#10 counter$count = 57028;
	#10 counter$count = 57029;
	#10 counter$count = 57030;
	#10 counter$count = 57031;
	#10 counter$count = 57032;
	#10 counter$count = 57033;
	#10 counter$count = 57034;
	#10 counter$count = 57035;
	#10 counter$count = 57036;
	#10 counter$count = 57037;
	#10 counter$count = 57038;
	#10 counter$count = 57039;
	#10 counter$count = 57040;
	#10 counter$count = 57041;
	#10 counter$count = 57042;
	#10 counter$count = 57043;
	#10 counter$count = 57044;
	#10 counter$count = 57045;
	#10 counter$count = 57046;
	#10 counter$count = 57047;
	#10 counter$count = 57048;
	#10 counter$count = 57049;
	#10 counter$count = 57050;
	#10 counter$count = 57051;
	#10 counter$count = 57052;
	#10 counter$count = 57053;
	#10 counter$count = 57054;
	#10 counter$count = 57055;
	#10 counter$count = 57056;
	#10 counter$count = 57057;
	#10 counter$count = 57058;
	#10 counter$count = 57059;
	#10 counter$count = 57060;
	#10 counter$count = 57061;
	#10 counter$count = 57062;
	#10 counter$count = 57063;
	#10 counter$count = 57064;
	#10 counter$count = 57065;
	#10 counter$count = 57066;
	#10 counter$count = 57067;
	#10 counter$count = 57068;
	#10 counter$count = 57069;
	#10 counter$count = 57070;
	#10 counter$count = 57071;
	#10 counter$count = 57072;
	#10 counter$count = 57073;
	#10 counter$count = 57074;
	#10 counter$count = 57075;
	#10 counter$count = 57076;
	#10 counter$count = 57077;
	#10 counter$count = 57078;
	#10 counter$count = 57079;
	#10 counter$count = 57080;
	#10 counter$count = 57081;
	#10 counter$count = 57082;
	#10 counter$count = 57083;
	#10 counter$count = 57084;
	#10 counter$count = 57085;
	#10 counter$count = 57086;
	#10 counter$count = 57087;
	#10 counter$count = 57088;
	#10 counter$count = 57089;
	#10 counter$count = 57090;
	#10 counter$count = 57091;
	#10 counter$count = 57092;
	#10 counter$count = 57093;
	#10 counter$count = 57094;
	#10 counter$count = 57095;
	#10 counter$count = 57096;
	#10 counter$count = 57097;
	#10 counter$count = 57098;
	#10 counter$count = 57099;
	#10 counter$count = 57100;
	#10 counter$count = 57101;
	#10 counter$count = 57102;
	#10 counter$count = 57103;
	#10 counter$count = 57104;
	#10 counter$count = 57105;
	#10 counter$count = 57106;
	#10 counter$count = 57107;
	#10 counter$count = 57108;
	#10 counter$count = 57109;
	#10 counter$count = 57110;
	#10 counter$count = 57111;
	#10 counter$count = 57112;
	#10 counter$count = 57113;
	#10 counter$count = 57114;
	#10 counter$count = 57115;
	#10 counter$count = 57116;
	#10 counter$count = 57117;
	#10 counter$count = 57118;
	#10 counter$count = 57119;
	#10 counter$count = 57120;
	#10 counter$count = 57121;
	#10 counter$count = 57122;
	#10 counter$count = 57123;
	#10 counter$count = 57124;
	#10 counter$count = 57125;
	#10 counter$count = 57126;
	#10 counter$count = 57127;
	#10 counter$count = 57128;
	#10 counter$count = 57129;
	#10 counter$count = 57130;
	#10 counter$count = 57131;
	#10 counter$count = 57132;
	#10 counter$count = 57133;
	#10 counter$count = 57134;
	#10 counter$count = 57135;
	#10 counter$count = 57136;
	#10 counter$count = 57137;
	#10 counter$count = 57138;
	#10 counter$count = 57139;
	#10 counter$count = 57140;
	#10 counter$count = 57141;
	#10 counter$count = 57142;
	#10 counter$count = 57143;
	#10 counter$count = 57144;
	#10 counter$count = 57145;
	#10 counter$count = 57146;
	#10 counter$count = 57147;
	#10 counter$count = 57148;
	#10 counter$count = 57149;
	#10 counter$count = 57150;
	#10 counter$count = 57151;
	#10 counter$count = 57152;
	#10 counter$count = 57153;
	#10 counter$count = 57154;
	#10 counter$count = 57155;
	#10 counter$count = 57156;
	#10 counter$count = 57157;
	#10 counter$count = 57158;
	#10 counter$count = 57159;
	#10 counter$count = 57160;
	#10 counter$count = 57161;
	#10 counter$count = 57162;
	#10 counter$count = 57163;
	#10 counter$count = 57164;
	#10 counter$count = 57165;
	#10 counter$count = 57166;
	#10 counter$count = 57167;
	#10 counter$count = 57168;
	#10 counter$count = 57169;
	#10 counter$count = 57170;
	#10 counter$count = 57171;
	#10 counter$count = 57172;
	#10 counter$count = 57173;
	#10 counter$count = 57174;
	#10 counter$count = 57175;
	#10 counter$count = 57176;
	#10 counter$count = 57177;
	#10 counter$count = 57178;
	#10 counter$count = 57179;
	#10 counter$count = 57180;
	#10 counter$count = 57181;
	#10 counter$count = 57182;
	#10 counter$count = 57183;
	#10 counter$count = 57184;
	#10 counter$count = 57185;
	#10 counter$count = 57186;
	#10 counter$count = 57187;
	#10 counter$count = 57188;
	#10 counter$count = 57189;
	#10 counter$count = 57190;
	#10 counter$count = 57191;
	#10 counter$count = 57192;
	#10 counter$count = 57193;
	#10 counter$count = 57194;
	#10 counter$count = 57195;
	#10 counter$count = 57196;
	#10 counter$count = 57197;
	#10 counter$count = 57198;
	#10 counter$count = 57199;
	#10 counter$count = 57200;
	#10 counter$count = 57201;
	#10 counter$count = 57202;
	#10 counter$count = 57203;
	#10 counter$count = 57204;
	#10 counter$count = 57205;
	#10 counter$count = 57206;
	#10 counter$count = 57207;
	#10 counter$count = 57208;
	#10 counter$count = 57209;
	#10 counter$count = 57210;
	#10 counter$count = 57211;
	#10 counter$count = 57212;
	#10 counter$count = 57213;
	#10 counter$count = 57214;
	#10 counter$count = 57215;
	#10 counter$count = 57216;
	#10 counter$count = 57217;
	#10 counter$count = 57218;
	#10 counter$count = 57219;
	#10 counter$count = 57220;
	#10 counter$count = 57221;
	#10 counter$count = 57222;
	#10 counter$count = 57223;
	#10 counter$count = 57224;
	#10 counter$count = 57225;
	#10 counter$count = 57226;
	#10 counter$count = 57227;
	#10 counter$count = 57228;
	#10 counter$count = 57229;
	#10 counter$count = 57230;
	#10 counter$count = 57231;
	#10 counter$count = 57232;
	#10 counter$count = 57233;
	#10 counter$count = 57234;
	#10 counter$count = 57235;
	#10 counter$count = 57236;
	#10 counter$count = 57237;
	#10 counter$count = 57238;
	#10 counter$count = 57239;
	#10 counter$count = 57240;
	#10 counter$count = 57241;
	#10 counter$count = 57242;
	#10 counter$count = 57243;
	#10 counter$count = 57244;
	#10 counter$count = 57245;
	#10 counter$count = 57246;
	#10 counter$count = 57247;
	#10 counter$count = 57248;
	#10 counter$count = 57249;
	#10 counter$count = 57250;
	#10 counter$count = 57251;
	#10 counter$count = 57252;
	#10 counter$count = 57253;
	#10 counter$count = 57254;
	#10 counter$count = 57255;
	#10 counter$count = 57256;
	#10 counter$count = 57257;
	#10 counter$count = 57258;
	#10 counter$count = 57259;
	#10 counter$count = 57260;
	#10 counter$count = 57261;
	#10 counter$count = 57262;
	#10 counter$count = 57263;
	#10 counter$count = 57264;
	#10 counter$count = 57265;
	#10 counter$count = 57266;
	#10 counter$count = 57267;
	#10 counter$count = 57268;
	#10 counter$count = 57269;
	#10 counter$count = 57270;
	#10 counter$count = 57271;
	#10 counter$count = 57272;
	#10 counter$count = 57273;
	#10 counter$count = 57274;
	#10 counter$count = 57275;
	#10 counter$count = 57276;
	#10 counter$count = 57277;
	#10 counter$count = 57278;
	#10 counter$count = 57279;
	#10 counter$count = 57280;
	#10 counter$count = 57281;
	#10 counter$count = 57282;
	#10 counter$count = 57283;
	#10 counter$count = 57284;
	#10 counter$count = 57285;
	#10 counter$count = 57286;
	#10 counter$count = 57287;
	#10 counter$count = 57288;
	#10 counter$count = 57289;
	#10 counter$count = 57290;
	#10 counter$count = 57291;
	#10 counter$count = 57292;
	#10 counter$count = 57293;
	#10 counter$count = 57294;
	#10 counter$count = 57295;
	#10 counter$count = 57296;
	#10 counter$count = 57297;
	#10 counter$count = 57298;
	#10 counter$count = 57299;
	#10 counter$count = 57300;
	#10 counter$count = 57301;
	#10 counter$count = 57302;
	#10 counter$count = 57303;
	#10 counter$count = 57304;
	#10 counter$count = 57305;
	#10 counter$count = 57306;
	#10 counter$count = 57307;
	#10 counter$count = 57308;
	#10 counter$count = 57309;
	#10 counter$count = 57310;
	#10 counter$count = 57311;
	#10 counter$count = 57312;
	#10 counter$count = 57313;
	#10 counter$count = 57314;
	#10 counter$count = 57315;
	#10 counter$count = 57316;
	#10 counter$count = 57317;
	#10 counter$count = 57318;
	#10 counter$count = 57319;
	#10 counter$count = 57320;
	#10 counter$count = 57321;
	#10 counter$count = 57322;
	#10 counter$count = 57323;
	#10 counter$count = 57324;
	#10 counter$count = 57325;
	#10 counter$count = 57326;
	#10 counter$count = 57327;
	#10 counter$count = 57328;
	#10 counter$count = 57329;
	#10 counter$count = 57330;
	#10 counter$count = 57331;
	#10 counter$count = 57332;
	#10 counter$count = 57333;
	#10 counter$count = 57334;
	#10 counter$count = 57335;
	#10 counter$count = 57336;
	#10 counter$count = 57337;
	#10 counter$count = 57338;
	#10 counter$count = 57339;
	#10 counter$count = 57340;
	#10 counter$count = 57341;
	#10 counter$count = 57342;
	#10 counter$count = 57343;
	#10 counter$count = 57344;
	#10 counter$count = 57345;
	#10 counter$count = 57346;
	#10 counter$count = 57347;
	#10 counter$count = 57348;
	#10 counter$count = 57349;
	#10 counter$count = 57350;
	#10 counter$count = 57351;
	#10 counter$count = 57352;
	#10 counter$count = 57353;
	#10 counter$count = 57354;
	#10 counter$count = 57355;
	#10 counter$count = 57356;
	#10 counter$count = 57357;
	#10 counter$count = 57358;
	#10 counter$count = 57359;
	#10 counter$count = 57360;
	#10 counter$count = 57361;
	#10 counter$count = 57362;
	#10 counter$count = 57363;
	#10 counter$count = 57364;
	#10 counter$count = 57365;
	#10 counter$count = 57366;
	#10 counter$count = 57367;
	#10 counter$count = 57368;
	#10 counter$count = 57369;
	#10 counter$count = 57370;
	#10 counter$count = 57371;
	#10 counter$count = 57372;
	#10 counter$count = 57373;
	#10 counter$count = 57374;
	#10 counter$count = 57375;
	#10 counter$count = 57376;
	#10 counter$count = 57377;
	#10 counter$count = 57378;
	#10 counter$count = 57379;
	#10 counter$count = 57380;
	#10 counter$count = 57381;
	#10 counter$count = 57382;
	#10 counter$count = 57383;
	#10 counter$count = 57384;
	#10 counter$count = 57385;
	#10 counter$count = 57386;
	#10 counter$count = 57387;
	#10 counter$count = 57388;
	#10 counter$count = 57389;
	#10 counter$count = 57390;
	#10 counter$count = 57391;
	#10 counter$count = 57392;
	#10 counter$count = 57393;
	#10 counter$count = 57394;
	#10 counter$count = 57395;
	#10 counter$count = 57396;
	#10 counter$count = 57397;
	#10 counter$count = 57398;
	#10 counter$count = 57399;
	#10 counter$count = 57400;
	#10 counter$count = 57401;
	#10 counter$count = 57402;
	#10 counter$count = 57403;
	#10 counter$count = 57404;
	#10 counter$count = 57405;
	#10 counter$count = 57406;
	#10 counter$count = 57407;
	#10 counter$count = 57408;
	#10 counter$count = 57409;
	#10 counter$count = 57410;
	#10 counter$count = 57411;
	#10 counter$count = 57412;
	#10 counter$count = 57413;
	#10 counter$count = 57414;
	#10 counter$count = 57415;
	#10 counter$count = 57416;
	#10 counter$count = 57417;
	#10 counter$count = 57418;
	#10 counter$count = 57419;
	#10 counter$count = 57420;
	#10 counter$count = 57421;
	#10 counter$count = 57422;
	#10 counter$count = 57423;
	#10 counter$count = 57424;
	#10 counter$count = 57425;
	#10 counter$count = 57426;
	#10 counter$count = 57427;
	#10 counter$count = 57428;
	#10 counter$count = 57429;
	#10 counter$count = 57430;
	#10 counter$count = 57431;
	#10 counter$count = 57432;
	#10 counter$count = 57433;
	#10 counter$count = 57434;
	#10 counter$count = 57435;
	#10 counter$count = 57436;
	#10 counter$count = 57437;
	#10 counter$count = 57438;
	#10 counter$count = 57439;
	#10 counter$count = 57440;
	#10 counter$count = 57441;
	#10 counter$count = 57442;
	#10 counter$count = 57443;
	#10 counter$count = 57444;
	#10 counter$count = 57445;
	#10 counter$count = 57446;
	#10 counter$count = 57447;
	#10 counter$count = 57448;
	#10 counter$count = 57449;
	#10 counter$count = 57450;
	#10 counter$count = 57451;
	#10 counter$count = 57452;
	#10 counter$count = 57453;
	#10 counter$count = 57454;
	#10 counter$count = 57455;
	#10 counter$count = 57456;
	#10 counter$count = 57457;
	#10 counter$count = 57458;
	#10 counter$count = 57459;
	#10 counter$count = 57460;
	#10 counter$count = 57461;
	#10 counter$count = 57462;
	#10 counter$count = 57463;
	#10 counter$count = 57464;
	#10 counter$count = 57465;
	#10 counter$count = 57466;
	#10 counter$count = 57467;
	#10 counter$count = 57468;
	#10 counter$count = 57469;
	#10 counter$count = 57470;
	#10 counter$count = 57471;
	#10 counter$count = 57472;
	#10 counter$count = 57473;
	#10 counter$count = 57474;
	#10 counter$count = 57475;
	#10 counter$count = 57476;
	#10 counter$count = 57477;
	#10 counter$count = 57478;
	#10 counter$count = 57479;
	#10 counter$count = 57480;
	#10 counter$count = 57481;
	#10 counter$count = 57482;
	#10 counter$count = 57483;
	#10 counter$count = 57484;
	#10 counter$count = 57485;
	#10 counter$count = 57486;
	#10 counter$count = 57487;
	#10 counter$count = 57488;
	#10 counter$count = 57489;
	#10 counter$count = 57490;
	#10 counter$count = 57491;
	#10 counter$count = 57492;
	#10 counter$count = 57493;
	#10 counter$count = 57494;
	#10 counter$count = 57495;
	#10 counter$count = 57496;
	#10 counter$count = 57497;
	#10 counter$count = 57498;
	#10 counter$count = 57499;
	#10 counter$count = 57500;
	#10 counter$count = 57501;
	#10 counter$count = 57502;
	#10 counter$count = 57503;
	#10 counter$count = 57504;
	#10 counter$count = 57505;
	#10 counter$count = 57506;
	#10 counter$count = 57507;
	#10 counter$count = 57508;
	#10 counter$count = 57509;
	#10 counter$count = 57510;
	#10 counter$count = 57511;
	#10 counter$count = 57512;
	#10 counter$count = 57513;
	#10 counter$count = 57514;
	#10 counter$count = 57515;
	#10 counter$count = 57516;
	#10 counter$count = 57517;
	#10 counter$count = 57518;
	#10 counter$count = 57519;
	#10 counter$count = 57520;
	#10 counter$count = 57521;
	#10 counter$count = 57522;
	#10 counter$count = 57523;
	#10 counter$count = 57524;
	#10 counter$count = 57525;
	#10 counter$count = 57526;
	#10 counter$count = 57527;
	#10 counter$count = 57528;
	#10 counter$count = 57529;
	#10 counter$count = 57530;
	#10 counter$count = 57531;
	#10 counter$count = 57532;
	#10 counter$count = 57533;
	#10 counter$count = 57534;
	#10 counter$count = 57535;
	#10 counter$count = 57536;
	#10 counter$count = 57537;
	#10 counter$count = 57538;
	#10 counter$count = 57539;
	#10 counter$count = 57540;
	#10 counter$count = 57541;
	#10 counter$count = 57542;
	#10 counter$count = 57543;
	#10 counter$count = 57544;
	#10 counter$count = 57545;
	#10 counter$count = 57546;
	#10 counter$count = 57547;
	#10 counter$count = 57548;
	#10 counter$count = 57549;
	#10 counter$count = 57550;
	#10 counter$count = 57551;
	#10 counter$count = 57552;
	#10 counter$count = 57553;
	#10 counter$count = 57554;
	#10 counter$count = 57555;
	#10 counter$count = 57556;
	#10 counter$count = 57557;
	#10 counter$count = 57558;
	#10 counter$count = 57559;
	#10 counter$count = 57560;
	#10 counter$count = 57561;
	#10 counter$count = 57562;
	#10 counter$count = 57563;
	#10 counter$count = 57564;
	#10 counter$count = 57565;
	#10 counter$count = 57566;
	#10 counter$count = 57567;
	#10 counter$count = 57568;
	#10 counter$count = 57569;
	#10 counter$count = 57570;
	#10 counter$count = 57571;
	#10 counter$count = 57572;
	#10 counter$count = 57573;
	#10 counter$count = 57574;
	#10 counter$count = 57575;
	#10 counter$count = 57576;
	#10 counter$count = 57577;
	#10 counter$count = 57578;
	#10 counter$count = 57579;
	#10 counter$count = 57580;
	#10 counter$count = 57581;
	#10 counter$count = 57582;
	#10 counter$count = 57583;
	#10 counter$count = 57584;
	#10 counter$count = 57585;
	#10 counter$count = 57586;
	#10 counter$count = 57587;
	#10 counter$count = 57588;
	#10 counter$count = 57589;
	#10 counter$count = 57590;
	#10 counter$count = 57591;
	#10 counter$count = 57592;
	#10 counter$count = 57593;
	#10 counter$count = 57594;
	#10 counter$count = 57595;
	#10 counter$count = 57596;
	#10 counter$count = 57597;
	#10 counter$count = 57598;
	#10 counter$count = 57599;
	#10 counter$count = 57600;
	#10 counter$count = 57601;
	#10 counter$count = 57602;
	#10 counter$count = 57603;
	#10 counter$count = 57604;
	#10 counter$count = 57605;
	#10 counter$count = 57606;
	#10 counter$count = 57607;
	#10 counter$count = 57608;
	#10 counter$count = 57609;
	#10 counter$count = 57610;
	#10 counter$count = 57611;
	#10 counter$count = 57612;
	#10 counter$count = 57613;
	#10 counter$count = 57614;
	#10 counter$count = 57615;
	#10 counter$count = 57616;
	#10 counter$count = 57617;
	#10 counter$count = 57618;
	#10 counter$count = 57619;
	#10 counter$count = 57620;
	#10 counter$count = 57621;
	#10 counter$count = 57622;
	#10 counter$count = 57623;
	#10 counter$count = 57624;
	#10 counter$count = 57625;
	#10 counter$count = 57626;
	#10 counter$count = 57627;
	#10 counter$count = 57628;
	#10 counter$count = 57629;
	#10 counter$count = 57630;
	#10 counter$count = 57631;
	#10 counter$count = 57632;
	#10 counter$count = 57633;
	#10 counter$count = 57634;
	#10 counter$count = 57635;
	#10 counter$count = 57636;
	#10 counter$count = 57637;
	#10 counter$count = 57638;
	#10 counter$count = 57639;
	#10 counter$count = 57640;
	#10 counter$count = 57641;
	#10 counter$count = 57642;
	#10 counter$count = 57643;
	#10 counter$count = 57644;
	#10 counter$count = 57645;
	#10 counter$count = 57646;
	#10 counter$count = 57647;
	#10 counter$count = 57648;
	#10 counter$count = 57649;
	#10 counter$count = 57650;
	#10 counter$count = 57651;
	#10 counter$count = 57652;
	#10 counter$count = 57653;
	#10 counter$count = 57654;
	#10 counter$count = 57655;
	#10 counter$count = 57656;
	#10 counter$count = 57657;
	#10 counter$count = 57658;
	#10 counter$count = 57659;
	#10 counter$count = 57660;
	#10 counter$count = 57661;
	#10 counter$count = 57662;
	#10 counter$count = 57663;
	#10 counter$count = 57664;
	#10 counter$count = 57665;
	#10 counter$count = 57666;
	#10 counter$count = 57667;
	#10 counter$count = 57668;
	#10 counter$count = 57669;
	#10 counter$count = 57670;
	#10 counter$count = 57671;
	#10 counter$count = 57672;
	#10 counter$count = 57673;
	#10 counter$count = 57674;
	#10 counter$count = 57675;
	#10 counter$count = 57676;
	#10 counter$count = 57677;
	#10 counter$count = 57678;
	#10 counter$count = 57679;
	#10 counter$count = 57680;
	#10 counter$count = 57681;
	#10 counter$count = 57682;
	#10 counter$count = 57683;
	#10 counter$count = 57684;
	#10 counter$count = 57685;
	#10 counter$count = 57686;
	#10 counter$count = 57687;
	#10 counter$count = 57688;
	#10 counter$count = 57689;
	#10 counter$count = 57690;
	#10 counter$count = 57691;
	#10 counter$count = 57692;
	#10 counter$count = 57693;
	#10 counter$count = 57694;
	#10 counter$count = 57695;
	#10 counter$count = 57696;
	#10 counter$count = 57697;
	#10 counter$count = 57698;
	#10 counter$count = 57699;
	#10 counter$count = 57700;
	#10 counter$count = 57701;
	#10 counter$count = 57702;
	#10 counter$count = 57703;
	#10 counter$count = 57704;
	#10 counter$count = 57705;
	#10 counter$count = 57706;
	#10 counter$count = 57707;
	#10 counter$count = 57708;
	#10 counter$count = 57709;
	#10 counter$count = 57710;
	#10 counter$count = 57711;
	#10 counter$count = 57712;
	#10 counter$count = 57713;
	#10 counter$count = 57714;
	#10 counter$count = 57715;
	#10 counter$count = 57716;
	#10 counter$count = 57717;
	#10 counter$count = 57718;
	#10 counter$count = 57719;
	#10 counter$count = 57720;
	#10 counter$count = 57721;
	#10 counter$count = 57722;
	#10 counter$count = 57723;
	#10 counter$count = 57724;
	#10 counter$count = 57725;
	#10 counter$count = 57726;
	#10 counter$count = 57727;
	#10 counter$count = 57728;
	#10 counter$count = 57729;
	#10 counter$count = 57730;
	#10 counter$count = 57731;
	#10 counter$count = 57732;
	#10 counter$count = 57733;
	#10 counter$count = 57734;
	#10 counter$count = 57735;
	#10 counter$count = 57736;
	#10 counter$count = 57737;
	#10 counter$count = 57738;
	#10 counter$count = 57739;
	#10 counter$count = 57740;
	#10 counter$count = 57741;
	#10 counter$count = 57742;
	#10 counter$count = 57743;
	#10 counter$count = 57744;
	#10 counter$count = 57745;
	#10 counter$count = 57746;
	#10 counter$count = 57747;
	#10 counter$count = 57748;
	#10 counter$count = 57749;
	#10 counter$count = 57750;
	#10 counter$count = 57751;
	#10 counter$count = 57752;
	#10 counter$count = 57753;
	#10 counter$count = 57754;
	#10 counter$count = 57755;
	#10 counter$count = 57756;
	#10 counter$count = 57757;
	#10 counter$count = 57758;
	#10 counter$count = 57759;
	#10 counter$count = 57760;
	#10 counter$count = 57761;
	#10 counter$count = 57762;
	#10 counter$count = 57763;
	#10 counter$count = 57764;
	#10 counter$count = 57765;
	#10 counter$count = 57766;
	#10 counter$count = 57767;
	#10 counter$count = 57768;
	#10 counter$count = 57769;
	#10 counter$count = 57770;
	#10 counter$count = 57771;
	#10 counter$count = 57772;
	#10 counter$count = 57773;
	#10 counter$count = 57774;
	#10 counter$count = 57775;
	#10 counter$count = 57776;
	#10 counter$count = 57777;
	#10 counter$count = 57778;
	#10 counter$count = 57779;
	#10 counter$count = 57780;
	#10 counter$count = 57781;
	#10 counter$count = 57782;
	#10 counter$count = 57783;
	#10 counter$count = 57784;
	#10 counter$count = 57785;
	#10 counter$count = 57786;
	#10 counter$count = 57787;
	#10 counter$count = 57788;
	#10 counter$count = 57789;
	#10 counter$count = 57790;
	#10 counter$count = 57791;
	#10 counter$count = 57792;
	#10 counter$count = 57793;
	#10 counter$count = 57794;
	#10 counter$count = 57795;
	#10 counter$count = 57796;
	#10 counter$count = 57797;
	#10 counter$count = 57798;
	#10 counter$count = 57799;
	#10 counter$count = 57800;
	#10 counter$count = 57801;
	#10 counter$count = 57802;
	#10 counter$count = 57803;
	#10 counter$count = 57804;
	#10 counter$count = 57805;
	#10 counter$count = 57806;
	#10 counter$count = 57807;
	#10 counter$count = 57808;
	#10 counter$count = 57809;
	#10 counter$count = 57810;
	#10 counter$count = 57811;
	#10 counter$count = 57812;
	#10 counter$count = 57813;
	#10 counter$count = 57814;
	#10 counter$count = 57815;
	#10 counter$count = 57816;
	#10 counter$count = 57817;
	#10 counter$count = 57818;
	#10 counter$count = 57819;
	#10 counter$count = 57820;
	#10 counter$count = 57821;
	#10 counter$count = 57822;
	#10 counter$count = 57823;
	#10 counter$count = 57824;
	#10 counter$count = 57825;
	#10 counter$count = 57826;
	#10 counter$count = 57827;
	#10 counter$count = 57828;
	#10 counter$count = 57829;
	#10 counter$count = 57830;
	#10 counter$count = 57831;
	#10 counter$count = 57832;
	#10 counter$count = 57833;
	#10 counter$count = 57834;
	#10 counter$count = 57835;
	#10 counter$count = 57836;
	#10 counter$count = 57837;
	#10 counter$count = 57838;
	#10 counter$count = 57839;
	#10 counter$count = 57840;
	#10 counter$count = 57841;
	#10 counter$count = 57842;
	#10 counter$count = 57843;
	#10 counter$count = 57844;
	#10 counter$count = 57845;
	#10 counter$count = 57846;
	#10 counter$count = 57847;
	#10 counter$count = 57848;
	#10 counter$count = 57849;
	#10 counter$count = 57850;
	#10 counter$count = 57851;
	#10 counter$count = 57852;
	#10 counter$count = 57853;
	#10 counter$count = 57854;
	#10 counter$count = 57855;
	#10 counter$count = 57856;
	#10 counter$count = 57857;
	#10 counter$count = 57858;
	#10 counter$count = 57859;
	#10 counter$count = 57860;
	#10 counter$count = 57861;
	#10 counter$count = 57862;
	#10 counter$count = 57863;
	#10 counter$count = 57864;
	#10 counter$count = 57865;
	#10 counter$count = 57866;
	#10 counter$count = 57867;
	#10 counter$count = 57868;
	#10 counter$count = 57869;
	#10 counter$count = 57870;
	#10 counter$count = 57871;
	#10 counter$count = 57872;
	#10 counter$count = 57873;
	#10 counter$count = 57874;
	#10 counter$count = 57875;
	#10 counter$count = 57876;
	#10 counter$count = 57877;
	#10 counter$count = 57878;
	#10 counter$count = 57879;
	#10 counter$count = 57880;
	#10 counter$count = 57881;
	#10 counter$count = 57882;
	#10 counter$count = 57883;
	#10 counter$count = 57884;
	#10 counter$count = 57885;
	#10 counter$count = 57886;
	#10 counter$count = 57887;
	#10 counter$count = 57888;
	#10 counter$count = 57889;
	#10 counter$count = 57890;
	#10 counter$count = 57891;
	#10 counter$count = 57892;
	#10 counter$count = 57893;
	#10 counter$count = 57894;
	#10 counter$count = 57895;
	#10 counter$count = 57896;
	#10 counter$count = 57897;
	#10 counter$count = 57898;
	#10 counter$count = 57899;
	#10 counter$count = 57900;
	#10 counter$count = 57901;
	#10 counter$count = 57902;
	#10 counter$count = 57903;
	#10 counter$count = 57904;
	#10 counter$count = 57905;
	#10 counter$count = 57906;
	#10 counter$count = 57907;
	#10 counter$count = 57908;
	#10 counter$count = 57909;
	#10 counter$count = 57910;
	#10 counter$count = 57911;
	#10 counter$count = 57912;
	#10 counter$count = 57913;
	#10 counter$count = 57914;
	#10 counter$count = 57915;
	#10 counter$count = 57916;
	#10 counter$count = 57917;
	#10 counter$count = 57918;
	#10 counter$count = 57919;
	#10 counter$count = 57920;
	#10 counter$count = 57921;
	#10 counter$count = 57922;
	#10 counter$count = 57923;
	#10 counter$count = 57924;
	#10 counter$count = 57925;
	#10 counter$count = 57926;
	#10 counter$count = 57927;
	#10 counter$count = 57928;
	#10 counter$count = 57929;
	#10 counter$count = 57930;
	#10 counter$count = 57931;
	#10 counter$count = 57932;
	#10 counter$count = 57933;
	#10 counter$count = 57934;
	#10 counter$count = 57935;
	#10 counter$count = 57936;
	#10 counter$count = 57937;
	#10 counter$count = 57938;
	#10 counter$count = 57939;
	#10 counter$count = 57940;
	#10 counter$count = 57941;
	#10 counter$count = 57942;
	#10 counter$count = 57943;
	#10 counter$count = 57944;
	#10 counter$count = 57945;
	#10 counter$count = 57946;
	#10 counter$count = 57947;
	#10 counter$count = 57948;
	#10 counter$count = 57949;
	#10 counter$count = 57950;
	#10 counter$count = 57951;
	#10 counter$count = 57952;
	#10 counter$count = 57953;
	#10 counter$count = 57954;
	#10 counter$count = 57955;
	#10 counter$count = 57956;
	#10 counter$count = 57957;
	#10 counter$count = 57958;
	#10 counter$count = 57959;
	#10 counter$count = 57960;
	#10 counter$count = 57961;
	#10 counter$count = 57962;
	#10 counter$count = 57963;
	#10 counter$count = 57964;
	#10 counter$count = 57965;
	#10 counter$count = 57966;
	#10 counter$count = 57967;
	#10 counter$count = 57968;
	#10 counter$count = 57969;
	#10 counter$count = 57970;
	#10 counter$count = 57971;
	#10 counter$count = 57972;
	#10 counter$count = 57973;
	#10 counter$count = 57974;
	#10 counter$count = 57975;
	#10 counter$count = 57976;
	#10 counter$count = 57977;
	#10 counter$count = 57978;
	#10 counter$count = 57979;
	#10 counter$count = 57980;
	#10 counter$count = 57981;
	#10 counter$count = 57982;
	#10 counter$count = 57983;
	#10 counter$count = 57984;
	#10 counter$count = 57985;
	#10 counter$count = 57986;
	#10 counter$count = 57987;
	#10 counter$count = 57988;
	#10 counter$count = 57989;
	#10 counter$count = 57990;
	#10 counter$count = 57991;
	#10 counter$count = 57992;
	#10 counter$count = 57993;
	#10 counter$count = 57994;
	#10 counter$count = 57995;
	#10 counter$count = 57996;
	#10 counter$count = 57997;
	#10 counter$count = 57998;
	#10 counter$count = 57999;
	#10 counter$count = 58000;
	#10 counter$count = 58001;
	#10 counter$count = 58002;
	#10 counter$count = 58003;
	#10 counter$count = 58004;
	#10 counter$count = 58005;
	#10 counter$count = 58006;
	#10 counter$count = 58007;
	#10 counter$count = 58008;
	#10 counter$count = 58009;
	#10 counter$count = 58010;
	#10 counter$count = 58011;
	#10 counter$count = 58012;
	#10 counter$count = 58013;
	#10 counter$count = 58014;
	#10 counter$count = 58015;
	#10 counter$count = 58016;
	#10 counter$count = 58017;
	#10 counter$count = 58018;
	#10 counter$count = 58019;
	#10 counter$count = 58020;
	#10 counter$count = 58021;
	#10 counter$count = 58022;
	#10 counter$count = 58023;
	#10 counter$count = 58024;
	#10 counter$count = 58025;
	#10 counter$count = 58026;
	#10 counter$count = 58027;
	#10 counter$count = 58028;
	#10 counter$count = 58029;
	#10 counter$count = 58030;
	#10 counter$count = 58031;
	#10 counter$count = 58032;
	#10 counter$count = 58033;
	#10 counter$count = 58034;
	#10 counter$count = 58035;
	#10 counter$count = 58036;
	#10 counter$count = 58037;
	#10 counter$count = 58038;
	#10 counter$count = 58039;
	#10 counter$count = 58040;
	#10 counter$count = 58041;
	#10 counter$count = 58042;
	#10 counter$count = 58043;
	#10 counter$count = 58044;
	#10 counter$count = 58045;
	#10 counter$count = 58046;
	#10 counter$count = 58047;
	#10 counter$count = 58048;
	#10 counter$count = 58049;
	#10 counter$count = 58050;
	#10 counter$count = 58051;
	#10 counter$count = 58052;
	#10 counter$count = 58053;
	#10 counter$count = 58054;
	#10 counter$count = 58055;
	#10 counter$count = 58056;
	#10 counter$count = 58057;
	#10 counter$count = 58058;
	#10 counter$count = 58059;
	#10 counter$count = 58060;
	#10 counter$count = 58061;
	#10 counter$count = 58062;
	#10 counter$count = 58063;
	#10 counter$count = 58064;
	#10 counter$count = 58065;
	#10 counter$count = 58066;
	#10 counter$count = 58067;
	#10 counter$count = 58068;
	#10 counter$count = 58069;
	#10 counter$count = 58070;
	#10 counter$count = 58071;
	#10 counter$count = 58072;
	#10 counter$count = 58073;
	#10 counter$count = 58074;
	#10 counter$count = 58075;
	#10 counter$count = 58076;
	#10 counter$count = 58077;
	#10 counter$count = 58078;
	#10 counter$count = 58079;
	#10 counter$count = 58080;
	#10 counter$count = 58081;
	#10 counter$count = 58082;
	#10 counter$count = 58083;
	#10 counter$count = 58084;
	#10 counter$count = 58085;
	#10 counter$count = 58086;
	#10 counter$count = 58087;
	#10 counter$count = 58088;
	#10 counter$count = 58089;
	#10 counter$count = 58090;
	#10 counter$count = 58091;
	#10 counter$count = 58092;
	#10 counter$count = 58093;
	#10 counter$count = 58094;
	#10 counter$count = 58095;
	#10 counter$count = 58096;
	#10 counter$count = 58097;
	#10 counter$count = 58098;
	#10 counter$count = 58099;
	#10 counter$count = 58100;
	#10 counter$count = 58101;
	#10 counter$count = 58102;
	#10 counter$count = 58103;
	#10 counter$count = 58104;
	#10 counter$count = 58105;
	#10 counter$count = 58106;
	#10 counter$count = 58107;
	#10 counter$count = 58108;
	#10 counter$count = 58109;
	#10 counter$count = 58110;
	#10 counter$count = 58111;
	#10 counter$count = 58112;
	#10 counter$count = 58113;
	#10 counter$count = 58114;
	#10 counter$count = 58115;
	#10 counter$count = 58116;
	#10 counter$count = 58117;
	#10 counter$count = 58118;
	#10 counter$count = 58119;
	#10 counter$count = 58120;
	#10 counter$count = 58121;
	#10 counter$count = 58122;
	#10 counter$count = 58123;
	#10 counter$count = 58124;
	#10 counter$count = 58125;
	#10 counter$count = 58126;
	#10 counter$count = 58127;
	#10 counter$count = 58128;
	#10 counter$count = 58129;
	#10 counter$count = 58130;
	#10 counter$count = 58131;
	#10 counter$count = 58132;
	#10 counter$count = 58133;
	#10 counter$count = 58134;
	#10 counter$count = 58135;
	#10 counter$count = 58136;
	#10 counter$count = 58137;
	#10 counter$count = 58138;
	#10 counter$count = 58139;
	#10 counter$count = 58140;
	#10 counter$count = 58141;
	#10 counter$count = 58142;
	#10 counter$count = 58143;
	#10 counter$count = 58144;
	#10 counter$count = 58145;
	#10 counter$count = 58146;
	#10 counter$count = 58147;
	#10 counter$count = 58148;
	#10 counter$count = 58149;
	#10 counter$count = 58150;
	#10 counter$count = 58151;
	#10 counter$count = 58152;
	#10 counter$count = 58153;
	#10 counter$count = 58154;
	#10 counter$count = 58155;
	#10 counter$count = 58156;
	#10 counter$count = 58157;
	#10 counter$count = 58158;
	#10 counter$count = 58159;
	#10 counter$count = 58160;
	#10 counter$count = 58161;
	#10 counter$count = 58162;
	#10 counter$count = 58163;
	#10 counter$count = 58164;
	#10 counter$count = 58165;
	#10 counter$count = 58166;
	#10 counter$count = 58167;
	#10 counter$count = 58168;
	#10 counter$count = 58169;
	#10 counter$count = 58170;
	#10 counter$count = 58171;
	#10 counter$count = 58172;
	#10 counter$count = 58173;
	#10 counter$count = 58174;
	#10 counter$count = 58175;
	#10 counter$count = 58176;
	#10 counter$count = 58177;
	#10 counter$count = 58178;
	#10 counter$count = 58179;
	#10 counter$count = 58180;
	#10 counter$count = 58181;
	#10 counter$count = 58182;
	#10 counter$count = 58183;
	#10 counter$count = 58184;
	#10 counter$count = 58185;
	#10 counter$count = 58186;
	#10 counter$count = 58187;
	#10 counter$count = 58188;
	#10 counter$count = 58189;
	#10 counter$count = 58190;
	#10 counter$count = 58191;
	#10 counter$count = 58192;
	#10 counter$count = 58193;
	#10 counter$count = 58194;
	#10 counter$count = 58195;
	#10 counter$count = 58196;
	#10 counter$count = 58197;
	#10 counter$count = 58198;
	#10 counter$count = 58199;
	#10 counter$count = 58200;
	#10 counter$count = 58201;
	#10 counter$count = 58202;
	#10 counter$count = 58203;
	#10 counter$count = 58204;
	#10 counter$count = 58205;
	#10 counter$count = 58206;
	#10 counter$count = 58207;
	#10 counter$count = 58208;
	#10 counter$count = 58209;
	#10 counter$count = 58210;
	#10 counter$count = 58211;
	#10 counter$count = 58212;
	#10 counter$count = 58213;
	#10 counter$count = 58214;
	#10 counter$count = 58215;
	#10 counter$count = 58216;
	#10 counter$count = 58217;
	#10 counter$count = 58218;
	#10 counter$count = 58219;
	#10 counter$count = 58220;
	#10 counter$count = 58221;
	#10 counter$count = 58222;
	#10 counter$count = 58223;
	#10 counter$count = 58224;
	#10 counter$count = 58225;
	#10 counter$count = 58226;
	#10 counter$count = 58227;
	#10 counter$count = 58228;
	#10 counter$count = 58229;
	#10 counter$count = 58230;
	#10 counter$count = 58231;
	#10 counter$count = 58232;
	#10 counter$count = 58233;
	#10 counter$count = 58234;
	#10 counter$count = 58235;
	#10 counter$count = 58236;
	#10 counter$count = 58237;
	#10 counter$count = 58238;
	#10 counter$count = 58239;
	#10 counter$count = 58240;
	#10 counter$count = 58241;
	#10 counter$count = 58242;
	#10 counter$count = 58243;
	#10 counter$count = 58244;
	#10 counter$count = 58245;
	#10 counter$count = 58246;
	#10 counter$count = 58247;
	#10 counter$count = 58248;
	#10 counter$count = 58249;
	#10 counter$count = 58250;
	#10 counter$count = 58251;
	#10 counter$count = 58252;
	#10 counter$count = 58253;
	#10 counter$count = 58254;
	#10 counter$count = 58255;
	#10 counter$count = 58256;
	#10 counter$count = 58257;
	#10 counter$count = 58258;
	#10 counter$count = 58259;
	#10 counter$count = 58260;
	#10 counter$count = 58261;
	#10 counter$count = 58262;
	#10 counter$count = 58263;
	#10 counter$count = 58264;
	#10 counter$count = 58265;
	#10 counter$count = 58266;
	#10 counter$count = 58267;
	#10 counter$count = 58268;
	#10 counter$count = 58269;
	#10 counter$count = 58270;
	#10 counter$count = 58271;
	#10 counter$count = 58272;
	#10 counter$count = 58273;
	#10 counter$count = 58274;
	#10 counter$count = 58275;
	#10 counter$count = 58276;
	#10 counter$count = 58277;
	#10 counter$count = 58278;
	#10 counter$count = 58279;
	#10 counter$count = 58280;
	#10 counter$count = 58281;
	#10 counter$count = 58282;
	#10 counter$count = 58283;
	#10 counter$count = 58284;
	#10 counter$count = 58285;
	#10 counter$count = 58286;
	#10 counter$count = 58287;
	#10 counter$count = 58288;
	#10 counter$count = 58289;
	#10 counter$count = 58290;
	#10 counter$count = 58291;
	#10 counter$count = 58292;
	#10 counter$count = 58293;
	#10 counter$count = 58294;
	#10 counter$count = 58295;
	#10 counter$count = 58296;
	#10 counter$count = 58297;
	#10 counter$count = 58298;
	#10 counter$count = 58299;
	#10 counter$count = 58300;
	#10 counter$count = 58301;
	#10 counter$count = 58302;
	#10 counter$count = 58303;
	#10 counter$count = 58304;
	#10 counter$count = 58305;
	#10 counter$count = 58306;
	#10 counter$count = 58307;
	#10 counter$count = 58308;
	#10 counter$count = 58309;
	#10 counter$count = 58310;
	#10 counter$count = 58311;
	#10 counter$count = 58312;
	#10 counter$count = 58313;
	#10 counter$count = 58314;
	#10 counter$count = 58315;
	#10 counter$count = 58316;
	#10 counter$count = 58317;
	#10 counter$count = 58318;
	#10 counter$count = 58319;
	#10 counter$count = 58320;
	#10 counter$count = 58321;
	#10 counter$count = 58322;
	#10 counter$count = 58323;
	#10 counter$count = 58324;
	#10 counter$count = 58325;
	#10 counter$count = 58326;
	#10 counter$count = 58327;
	#10 counter$count = 58328;
	#10 counter$count = 58329;
	#10 counter$count = 58330;
	#10 counter$count = 58331;
	#10 counter$count = 58332;
	#10 counter$count = 58333;
	#10 counter$count = 58334;
	#10 counter$count = 58335;
	#10 counter$count = 58336;
	#10 counter$count = 58337;
	#10 counter$count = 58338;
	#10 counter$count = 58339;
	#10 counter$count = 58340;
	#10 counter$count = 58341;
	#10 counter$count = 58342;
	#10 counter$count = 58343;
	#10 counter$count = 58344;
	#10 counter$count = 58345;
	#10 counter$count = 58346;
	#10 counter$count = 58347;
	#10 counter$count = 58348;
	#10 counter$count = 58349;
	#10 counter$count = 58350;
	#10 counter$count = 58351;
	#10 counter$count = 58352;
	#10 counter$count = 58353;
	#10 counter$count = 58354;
	#10 counter$count = 58355;
	#10 counter$count = 58356;
	#10 counter$count = 58357;
	#10 counter$count = 58358;
	#10 counter$count = 58359;
	#10 counter$count = 58360;
	#10 counter$count = 58361;
	#10 counter$count = 58362;
	#10 counter$count = 58363;
	#10 counter$count = 58364;
	#10 counter$count = 58365;
	#10 counter$count = 58366;
	#10 counter$count = 58367;
	#10 counter$count = 58368;
	#10 counter$count = 58369;
	#10 counter$count = 58370;
	#10 counter$count = 58371;
	#10 counter$count = 58372;
	#10 counter$count = 58373;
	#10 counter$count = 58374;
	#10 counter$count = 58375;
	#10 counter$count = 58376;
	#10 counter$count = 58377;
	#10 counter$count = 58378;
	#10 counter$count = 58379;
	#10 counter$count = 58380;
	#10 counter$count = 58381;
	#10 counter$count = 58382;
	#10 counter$count = 58383;
	#10 counter$count = 58384;
	#10 counter$count = 58385;
	#10 counter$count = 58386;
	#10 counter$count = 58387;
	#10 counter$count = 58388;
	#10 counter$count = 58389;
	#10 counter$count = 58390;
	#10 counter$count = 58391;
	#10 counter$count = 58392;
	#10 counter$count = 58393;
	#10 counter$count = 58394;
	#10 counter$count = 58395;
	#10 counter$count = 58396;
	#10 counter$count = 58397;
	#10 counter$count = 58398;
	#10 counter$count = 58399;
	#10 counter$count = 58400;
	#10 counter$count = 58401;
	#10 counter$count = 58402;
	#10 counter$count = 58403;
	#10 counter$count = 58404;
	#10 counter$count = 58405;
	#10 counter$count = 58406;
	#10 counter$count = 58407;
	#10 counter$count = 58408;
	#10 counter$count = 58409;
	#10 counter$count = 58410;
	#10 counter$count = 58411;
	#10 counter$count = 58412;
	#10 counter$count = 58413;
	#10 counter$count = 58414;
	#10 counter$count = 58415;
	#10 counter$count = 58416;
	#10 counter$count = 58417;
	#10 counter$count = 58418;
	#10 counter$count = 58419;
	#10 counter$count = 58420;
	#10 counter$count = 58421;
	#10 counter$count = 58422;
	#10 counter$count = 58423;
	#10 counter$count = 58424;
	#10 counter$count = 58425;
	#10 counter$count = 58426;
	#10 counter$count = 58427;
	#10 counter$count = 58428;
	#10 counter$count = 58429;
	#10 counter$count = 58430;
	#10 counter$count = 58431;
	#10 counter$count = 58432;
	#10 counter$count = 58433;
	#10 counter$count = 58434;
	#10 counter$count = 58435;
	#10 counter$count = 58436;
	#10 counter$count = 58437;
	#10 counter$count = 58438;
	#10 counter$count = 58439;
	#10 counter$count = 58440;
	#10 counter$count = 58441;
	#10 counter$count = 58442;
	#10 counter$count = 58443;
	#10 counter$count = 58444;
	#10 counter$count = 58445;
	#10 counter$count = 58446;
	#10 counter$count = 58447;
	#10 counter$count = 58448;
	#10 counter$count = 58449;
	#10 counter$count = 58450;
	#10 counter$count = 58451;
	#10 counter$count = 58452;
	#10 counter$count = 58453;
	#10 counter$count = 58454;
	#10 counter$count = 58455;
	#10 counter$count = 58456;
	#10 counter$count = 58457;
	#10 counter$count = 58458;
	#10 counter$count = 58459;
	#10 counter$count = 58460;
	#10 counter$count = 58461;
	#10 counter$count = 58462;
	#10 counter$count = 58463;
	#10 counter$count = 58464;
	#10 counter$count = 58465;
	#10 counter$count = 58466;
	#10 counter$count = 58467;
	#10 counter$count = 58468;
	#10 counter$count = 58469;
	#10 counter$count = 58470;
	#10 counter$count = 58471;
	#10 counter$count = 58472;
	#10 counter$count = 58473;
	#10 counter$count = 58474;
	#10 counter$count = 58475;
	#10 counter$count = 58476;
	#10 counter$count = 58477;
	#10 counter$count = 58478;
	#10 counter$count = 58479;
	#10 counter$count = 58480;
	#10 counter$count = 58481;
	#10 counter$count = 58482;
	#10 counter$count = 58483;
	#10 counter$count = 58484;
	#10 counter$count = 58485;
	#10 counter$count = 58486;
	#10 counter$count = 58487;
	#10 counter$count = 58488;
	#10 counter$count = 58489;
	#10 counter$count = 58490;
	#10 counter$count = 58491;
	#10 counter$count = 58492;
	#10 counter$count = 58493;
	#10 counter$count = 58494;
	#10 counter$count = 58495;
	#10 counter$count = 58496;
	#10 counter$count = 58497;
	#10 counter$count = 58498;
	#10 counter$count = 58499;
	#10 counter$count = 58500;
	#10 counter$count = 58501;
	#10 counter$count = 58502;
	#10 counter$count = 58503;
	#10 counter$count = 58504;
	#10 counter$count = 58505;
	#10 counter$count = 58506;
	#10 counter$count = 58507;
	#10 counter$count = 58508;
	#10 counter$count = 58509;
	#10 counter$count = 58510;
	#10 counter$count = 58511;
	#10 counter$count = 58512;
	#10 counter$count = 58513;
	#10 counter$count = 58514;
	#10 counter$count = 58515;
	#10 counter$count = 58516;
	#10 counter$count = 58517;
	#10 counter$count = 58518;
	#10 counter$count = 58519;
	#10 counter$count = 58520;
	#10 counter$count = 58521;
	#10 counter$count = 58522;
	#10 counter$count = 58523;
	#10 counter$count = 58524;
	#10 counter$count = 58525;
	#10 counter$count = 58526;
	#10 counter$count = 58527;
	#10 counter$count = 58528;
	#10 counter$count = 58529;
	#10 counter$count = 58530;
	#10 counter$count = 58531;
	#10 counter$count = 58532;
	#10 counter$count = 58533;
	#10 counter$count = 58534;
	#10 counter$count = 58535;
	#10 counter$count = 58536;
	#10 counter$count = 58537;
	#10 counter$count = 58538;
	#10 counter$count = 58539;
	#10 counter$count = 58540;
	#10 counter$count = 58541;
	#10 counter$count = 58542;
	#10 counter$count = 58543;
	#10 counter$count = 58544;
	#10 counter$count = 58545;
	#10 counter$count = 58546;
	#10 counter$count = 58547;
	#10 counter$count = 58548;
	#10 counter$count = 58549;
	#10 counter$count = 58550;
	#10 counter$count = 58551;
	#10 counter$count = 58552;
	#10 counter$count = 58553;
	#10 counter$count = 58554;
	#10 counter$count = 58555;
	#10 counter$count = 58556;
	#10 counter$count = 58557;
	#10 counter$count = 58558;
	#10 counter$count = 58559;
	#10 counter$count = 58560;
	#10 counter$count = 58561;
	#10 counter$count = 58562;
	#10 counter$count = 58563;
	#10 counter$count = 58564;
	#10 counter$count = 58565;
	#10 counter$count = 58566;
	#10 counter$count = 58567;
	#10 counter$count = 58568;
	#10 counter$count = 58569;
	#10 counter$count = 58570;
	#10 counter$count = 58571;
	#10 counter$count = 58572;
	#10 counter$count = 58573;
	#10 counter$count = 58574;
	#10 counter$count = 58575;
	#10 counter$count = 58576;
	#10 counter$count = 58577;
	#10 counter$count = 58578;
	#10 counter$count = 58579;
	#10 counter$count = 58580;
	#10 counter$count = 58581;
	#10 counter$count = 58582;
	#10 counter$count = 58583;
	#10 counter$count = 58584;
	#10 counter$count = 58585;
	#10 counter$count = 58586;
	#10 counter$count = 58587;
	#10 counter$count = 58588;
	#10 counter$count = 58589;
	#10 counter$count = 58590;
	#10 counter$count = 58591;
	#10 counter$count = 58592;
	#10 counter$count = 58593;
	#10 counter$count = 58594;
	#10 counter$count = 58595;
	#10 counter$count = 58596;
	#10 counter$count = 58597;
	#10 counter$count = 58598;
	#10 counter$count = 58599;
	#10 counter$count = 58600;
	#10 counter$count = 58601;
	#10 counter$count = 58602;
	#10 counter$count = 58603;
	#10 counter$count = 58604;
	#10 counter$count = 58605;
	#10 counter$count = 58606;
	#10 counter$count = 58607;
	#10 counter$count = 58608;
	#10 counter$count = 58609;
	#10 counter$count = 58610;
	#10 counter$count = 58611;
	#10 counter$count = 58612;
	#10 counter$count = 58613;
	#10 counter$count = 58614;
	#10 counter$count = 58615;
	#10 counter$count = 58616;
	#10 counter$count = 58617;
	#10 counter$count = 58618;
	#10 counter$count = 58619;
	#10 counter$count = 58620;
	#10 counter$count = 58621;
	#10 counter$count = 58622;
	#10 counter$count = 58623;
	#10 counter$count = 58624;
	#10 counter$count = 58625;
	#10 counter$count = 58626;
	#10 counter$count = 58627;
	#10 counter$count = 58628;
	#10 counter$count = 58629;
	#10 counter$count = 58630;
	#10 counter$count = 58631;
	#10 counter$count = 58632;
	#10 counter$count = 58633;
	#10 counter$count = 58634;
	#10 counter$count = 58635;
	#10 counter$count = 58636;
	#10 counter$count = 58637;
	#10 counter$count = 58638;
	#10 counter$count = 58639;
	#10 counter$count = 58640;
	#10 counter$count = 58641;
	#10 counter$count = 58642;
	#10 counter$count = 58643;
	#10 counter$count = 58644;
	#10 counter$count = 58645;
	#10 counter$count = 58646;
	#10 counter$count = 58647;
	#10 counter$count = 58648;
	#10 counter$count = 58649;
	#10 counter$count = 58650;
	#10 counter$count = 58651;
	#10 counter$count = 58652;
	#10 counter$count = 58653;
	#10 counter$count = 58654;
	#10 counter$count = 58655;
	#10 counter$count = 58656;
	#10 counter$count = 58657;
	#10 counter$count = 58658;
	#10 counter$count = 58659;
	#10 counter$count = 58660;
	#10 counter$count = 58661;
	#10 counter$count = 58662;
	#10 counter$count = 58663;
	#10 counter$count = 58664;
	#10 counter$count = 58665;
	#10 counter$count = 58666;
	#10 counter$count = 58667;
	#10 counter$count = 58668;
	#10 counter$count = 58669;
	#10 counter$count = 58670;
	#10 counter$count = 58671;
	#10 counter$count = 58672;
	#10 counter$count = 58673;
	#10 counter$count = 58674;
	#10 counter$count = 58675;
	#10 counter$count = 58676;
	#10 counter$count = 58677;
	#10 counter$count = 58678;
	#10 counter$count = 58679;
	#10 counter$count = 58680;
	#10 counter$count = 58681;
	#10 counter$count = 58682;
	#10 counter$count = 58683;
	#10 counter$count = 58684;
	#10 counter$count = 58685;
	#10 counter$count = 58686;
	#10 counter$count = 58687;
	#10 counter$count = 58688;
	#10 counter$count = 58689;
	#10 counter$count = 58690;
	#10 counter$count = 58691;
	#10 counter$count = 58692;
	#10 counter$count = 58693;
	#10 counter$count = 58694;
	#10 counter$count = 58695;
	#10 counter$count = 58696;
	#10 counter$count = 58697;
	#10 counter$count = 58698;
	#10 counter$count = 58699;
	#10 counter$count = 58700;
	#10 counter$count = 58701;
	#10 counter$count = 58702;
	#10 counter$count = 58703;
	#10 counter$count = 58704;
	#10 counter$count = 58705;
	#10 counter$count = 58706;
	#10 counter$count = 58707;
	#10 counter$count = 58708;
	#10 counter$count = 58709;
	#10 counter$count = 58710;
	#10 counter$count = 58711;
	#10 counter$count = 58712;
	#10 counter$count = 58713;
	#10 counter$count = 58714;
	#10 counter$count = 58715;
	#10 counter$count = 58716;
	#10 counter$count = 58717;
	#10 counter$count = 58718;
	#10 counter$count = 58719;
	#10 counter$count = 58720;
	#10 counter$count = 58721;
	#10 counter$count = 58722;
	#10 counter$count = 58723;
	#10 counter$count = 58724;
	#10 counter$count = 58725;
	#10 counter$count = 58726;
	#10 counter$count = 58727;
	#10 counter$count = 58728;
	#10 counter$count = 58729;
	#10 counter$count = 58730;
	#10 counter$count = 58731;
	#10 counter$count = 58732;
	#10 counter$count = 58733;
	#10 counter$count = 58734;
	#10 counter$count = 58735;
	#10 counter$count = 58736;
	#10 counter$count = 58737;
	#10 counter$count = 58738;
	#10 counter$count = 58739;
	#10 counter$count = 58740;
	#10 counter$count = 58741;
	#10 counter$count = 58742;
	#10 counter$count = 58743;
	#10 counter$count = 58744;
	#10 counter$count = 58745;
	#10 counter$count = 58746;
	#10 counter$count = 58747;
	#10 counter$count = 58748;
	#10 counter$count = 58749;
	#10 counter$count = 58750;
	#10 counter$count = 58751;
	#10 counter$count = 58752;
	#10 counter$count = 58753;
	#10 counter$count = 58754;
	#10 counter$count = 58755;
	#10 counter$count = 58756;
	#10 counter$count = 58757;
	#10 counter$count = 58758;
	#10 counter$count = 58759;
	#10 counter$count = 58760;
	#10 counter$count = 58761;
	#10 counter$count = 58762;
	#10 counter$count = 58763;
	#10 counter$count = 58764;
	#10 counter$count = 58765;
	#10 counter$count = 58766;
	#10 counter$count = 58767;
	#10 counter$count = 58768;
	#10 counter$count = 58769;
	#10 counter$count = 58770;
	#10 counter$count = 58771;
	#10 counter$count = 58772;
	#10 counter$count = 58773;
	#10 counter$count = 58774;
	#10 counter$count = 58775;
	#10 counter$count = 58776;
	#10 counter$count = 58777;
	#10 counter$count = 58778;
	#10 counter$count = 58779;
	#10 counter$count = 58780;
	#10 counter$count = 58781;
	#10 counter$count = 58782;
	#10 counter$count = 58783;
	#10 counter$count = 58784;
	#10 counter$count = 58785;
	#10 counter$count = 58786;
	#10 counter$count = 58787;
	#10 counter$count = 58788;
	#10 counter$count = 58789;
	#10 counter$count = 58790;
	#10 counter$count = 58791;
	#10 counter$count = 58792;
	#10 counter$count = 58793;
	#10 counter$count = 58794;
	#10 counter$count = 58795;
	#10 counter$count = 58796;
	#10 counter$count = 58797;
	#10 counter$count = 58798;
	#10 counter$count = 58799;
	#10 counter$count = 58800;
	#10 counter$count = 58801;
	#10 counter$count = 58802;
	#10 counter$count = 58803;
	#10 counter$count = 58804;
	#10 counter$count = 58805;
	#10 counter$count = 58806;
	#10 counter$count = 58807;
	#10 counter$count = 58808;
	#10 counter$count = 58809;
	#10 counter$count = 58810;
	#10 counter$count = 58811;
	#10 counter$count = 58812;
	#10 counter$count = 58813;
	#10 counter$count = 58814;
	#10 counter$count = 58815;
	#10 counter$count = 58816;
	#10 counter$count = 58817;
	#10 counter$count = 58818;
	#10 counter$count = 58819;
	#10 counter$count = 58820;
	#10 counter$count = 58821;
	#10 counter$count = 58822;
	#10 counter$count = 58823;
	#10 counter$count = 58824;
	#10 counter$count = 58825;
	#10 counter$count = 58826;
	#10 counter$count = 58827;
	#10 counter$count = 58828;
	#10 counter$count = 58829;
	#10 counter$count = 58830;
	#10 counter$count = 58831;
	#10 counter$count = 58832;
	#10 counter$count = 58833;
	#10 counter$count = 58834;
	#10 counter$count = 58835;
	#10 counter$count = 58836;
	#10 counter$count = 58837;
	#10 counter$count = 58838;
	#10 counter$count = 58839;
	#10 counter$count = 58840;
	#10 counter$count = 58841;
	#10 counter$count = 58842;
	#10 counter$count = 58843;
	#10 counter$count = 58844;
	#10 counter$count = 58845;
	#10 counter$count = 58846;
	#10 counter$count = 58847;
	#10 counter$count = 58848;
	#10 counter$count = 58849;
	#10 counter$count = 58850;
	#10 counter$count = 58851;
	#10 counter$count = 58852;
	#10 counter$count = 58853;
	#10 counter$count = 58854;
	#10 counter$count = 58855;
	#10 counter$count = 58856;
	#10 counter$count = 58857;
	#10 counter$count = 58858;
	#10 counter$count = 58859;
	#10 counter$count = 58860;
	#10 counter$count = 58861;
	#10 counter$count = 58862;
	#10 counter$count = 58863;
	#10 counter$count = 58864;
	#10 counter$count = 58865;
	#10 counter$count = 58866;
	#10 counter$count = 58867;
	#10 counter$count = 58868;
	#10 counter$count = 58869;
	#10 counter$count = 58870;
	#10 counter$count = 58871;
	#10 counter$count = 58872;
	#10 counter$count = 58873;
	#10 counter$count = 58874;
	#10 counter$count = 58875;
	#10 counter$count = 58876;
	#10 counter$count = 58877;
	#10 counter$count = 58878;
	#10 counter$count = 58879;
	#10 counter$count = 58880;
	#10 counter$count = 58881;
	#10 counter$count = 58882;
	#10 counter$count = 58883;
	#10 counter$count = 58884;
	#10 counter$count = 58885;
	#10 counter$count = 58886;
	#10 counter$count = 58887;
	#10 counter$count = 58888;
	#10 counter$count = 58889;
	#10 counter$count = 58890;
	#10 counter$count = 58891;
	#10 counter$count = 58892;
	#10 counter$count = 58893;
	#10 counter$count = 58894;
	#10 counter$count = 58895;
	#10 counter$count = 58896;
	#10 counter$count = 58897;
	#10 counter$count = 58898;
	#10 counter$count = 58899;
	#10 counter$count = 58900;
	#10 counter$count = 58901;
	#10 counter$count = 58902;
	#10 counter$count = 58903;
	#10 counter$count = 58904;
	#10 counter$count = 58905;
	#10 counter$count = 58906;
	#10 counter$count = 58907;
	#10 counter$count = 58908;
	#10 counter$count = 58909;
	#10 counter$count = 58910;
	#10 counter$count = 58911;
	#10 counter$count = 58912;
	#10 counter$count = 58913;
	#10 counter$count = 58914;
	#10 counter$count = 58915;
	#10 counter$count = 58916;
	#10 counter$count = 58917;
	#10 counter$count = 58918;
	#10 counter$count = 58919;
	#10 counter$count = 58920;
	#10 counter$count = 58921;
	#10 counter$count = 58922;
	#10 counter$count = 58923;
	#10 counter$count = 58924;
	#10 counter$count = 58925;
	#10 counter$count = 58926;
	#10 counter$count = 58927;
	#10 counter$count = 58928;
	#10 counter$count = 58929;
	#10 counter$count = 58930;
	#10 counter$count = 58931;
	#10 counter$count = 58932;
	#10 counter$count = 58933;
	#10 counter$count = 58934;
	#10 counter$count = 58935;
	#10 counter$count = 58936;
	#10 counter$count = 58937;
	#10 counter$count = 58938;
	#10 counter$count = 58939;
	#10 counter$count = 58940;
	#10 counter$count = 58941;
	#10 counter$count = 58942;
	#10 counter$count = 58943;
	#10 counter$count = 58944;
	#10 counter$count = 58945;
	#10 counter$count = 58946;
	#10 counter$count = 58947;
	#10 counter$count = 58948;
	#10 counter$count = 58949;
	#10 counter$count = 58950;
	#10 counter$count = 58951;
	#10 counter$count = 58952;
	#10 counter$count = 58953;
	#10 counter$count = 58954;
	#10 counter$count = 58955;
	#10 counter$count = 58956;
	#10 counter$count = 58957;
	#10 counter$count = 58958;
	#10 counter$count = 58959;
	#10 counter$count = 58960;
	#10 counter$count = 58961;
	#10 counter$count = 58962;
	#10 counter$count = 58963;
	#10 counter$count = 58964;
	#10 counter$count = 58965;
	#10 counter$count = 58966;
	#10 counter$count = 58967;
	#10 counter$count = 58968;
	#10 counter$count = 58969;
	#10 counter$count = 58970;
	#10 counter$count = 58971;
	#10 counter$count = 58972;
	#10 counter$count = 58973;
	#10 counter$count = 58974;
	#10 counter$count = 58975;
	#10 counter$count = 58976;
	#10 counter$count = 58977;
	#10 counter$count = 58978;
	#10 counter$count = 58979;
	#10 counter$count = 58980;
	#10 counter$count = 58981;
	#10 counter$count = 58982;
	#10 counter$count = 58983;
	#10 counter$count = 58984;
	#10 counter$count = 58985;
	#10 counter$count = 58986;
	#10 counter$count = 58987;
	#10 counter$count = 58988;
	#10 counter$count = 58989;
	#10 counter$count = 58990;
	#10 counter$count = 58991;
	#10 counter$count = 58992;
	#10 counter$count = 58993;
	#10 counter$count = 58994;
	#10 counter$count = 58995;
	#10 counter$count = 58996;
	#10 counter$count = 58997;
	#10 counter$count = 58998;
	#10 counter$count = 58999;
	#10 counter$count = 59000;
	#10 counter$count = 59001;
	#10 counter$count = 59002;
	#10 counter$count = 59003;
	#10 counter$count = 59004;
	#10 counter$count = 59005;
	#10 counter$count = 59006;
	#10 counter$count = 59007;
	#10 counter$count = 59008;
	#10 counter$count = 59009;
	#10 counter$count = 59010;
	#10 counter$count = 59011;
	#10 counter$count = 59012;
	#10 counter$count = 59013;
	#10 counter$count = 59014;
	#10 counter$count = 59015;
	#10 counter$count = 59016;
	#10 counter$count = 59017;
	#10 counter$count = 59018;
	#10 counter$count = 59019;
	#10 counter$count = 59020;
	#10 counter$count = 59021;
	#10 counter$count = 59022;
	#10 counter$count = 59023;
	#10 counter$count = 59024;
	#10 counter$count = 59025;
	#10 counter$count = 59026;
	#10 counter$count = 59027;
	#10 counter$count = 59028;
	#10 counter$count = 59029;
	#10 counter$count = 59030;
	#10 counter$count = 59031;
	#10 counter$count = 59032;
	#10 counter$count = 59033;
	#10 counter$count = 59034;
	#10 counter$count = 59035;
	#10 counter$count = 59036;
	#10 counter$count = 59037;
	#10 counter$count = 59038;
	#10 counter$count = 59039;
	#10 counter$count = 59040;
	#10 counter$count = 59041;
	#10 counter$count = 59042;
	#10 counter$count = 59043;
	#10 counter$count = 59044;
	#10 counter$count = 59045;
	#10 counter$count = 59046;
	#10 counter$count = 59047;
	#10 counter$count = 59048;
	#10 counter$count = 59049;
	#10 counter$count = 59050;
	#10 counter$count = 59051;
	#10 counter$count = 59052;
	#10 counter$count = 59053;
	#10 counter$count = 59054;
	#10 counter$count = 59055;
	#10 counter$count = 59056;
	#10 counter$count = 59057;
	#10 counter$count = 59058;
	#10 counter$count = 59059;
	#10 counter$count = 59060;
	#10 counter$count = 59061;
	#10 counter$count = 59062;
	#10 counter$count = 59063;
	#10 counter$count = 59064;
	#10 counter$count = 59065;
	#10 counter$count = 59066;
	#10 counter$count = 59067;
	#10 counter$count = 59068;
	#10 counter$count = 59069;
	#10 counter$count = 59070;
	#10 counter$count = 59071;
	#10 counter$count = 59072;
	#10 counter$count = 59073;
	#10 counter$count = 59074;
	#10 counter$count = 59075;
	#10 counter$count = 59076;
	#10 counter$count = 59077;
	#10 counter$count = 59078;
	#10 counter$count = 59079;
	#10 counter$count = 59080;
	#10 counter$count = 59081;
	#10 counter$count = 59082;
	#10 counter$count = 59083;
	#10 counter$count = 59084;
	#10 counter$count = 59085;
	#10 counter$count = 59086;
	#10 counter$count = 59087;
	#10 counter$count = 59088;
	#10 counter$count = 59089;
	#10 counter$count = 59090;
	#10 counter$count = 59091;
	#10 counter$count = 59092;
	#10 counter$count = 59093;
	#10 counter$count = 59094;
	#10 counter$count = 59095;
	#10 counter$count = 59096;
	#10 counter$count = 59097;
	#10 counter$count = 59098;
	#10 counter$count = 59099;
	#10 counter$count = 59100;
	#10 counter$count = 59101;
	#10 counter$count = 59102;
	#10 counter$count = 59103;
	#10 counter$count = 59104;
	#10 counter$count = 59105;
	#10 counter$count = 59106;
	#10 counter$count = 59107;
	#10 counter$count = 59108;
	#10 counter$count = 59109;
	#10 counter$count = 59110;
	#10 counter$count = 59111;
	#10 counter$count = 59112;
	#10 counter$count = 59113;
	#10 counter$count = 59114;
	#10 counter$count = 59115;
	#10 counter$count = 59116;
	#10 counter$count = 59117;
	#10 counter$count = 59118;
	#10 counter$count = 59119;
	#10 counter$count = 59120;
	#10 counter$count = 59121;
	#10 counter$count = 59122;
	#10 counter$count = 59123;
	#10 counter$count = 59124;
	#10 counter$count = 59125;
	#10 counter$count = 59126;
	#10 counter$count = 59127;
	#10 counter$count = 59128;
	#10 counter$count = 59129;
	#10 counter$count = 59130;
	#10 counter$count = 59131;
	#10 counter$count = 59132;
	#10 counter$count = 59133;
	#10 counter$count = 59134;
	#10 counter$count = 59135;
	#10 counter$count = 59136;
	#10 counter$count = 59137;
	#10 counter$count = 59138;
	#10 counter$count = 59139;
	#10 counter$count = 59140;
	#10 counter$count = 59141;
	#10 counter$count = 59142;
	#10 counter$count = 59143;
	#10 counter$count = 59144;
	#10 counter$count = 59145;
	#10 counter$count = 59146;
	#10 counter$count = 59147;
	#10 counter$count = 59148;
	#10 counter$count = 59149;
	#10 counter$count = 59150;
	#10 counter$count = 59151;
	#10 counter$count = 59152;
	#10 counter$count = 59153;
	#10 counter$count = 59154;
	#10 counter$count = 59155;
	#10 counter$count = 59156;
	#10 counter$count = 59157;
	#10 counter$count = 59158;
	#10 counter$count = 59159;
	#10 counter$count = 59160;
	#10 counter$count = 59161;
	#10 counter$count = 59162;
	#10 counter$count = 59163;
	#10 counter$count = 59164;
	#10 counter$count = 59165;
	#10 counter$count = 59166;
	#10 counter$count = 59167;
	#10 counter$count = 59168;
	#10 counter$count = 59169;
	#10 counter$count = 59170;
	#10 counter$count = 59171;
	#10 counter$count = 59172;
	#10 counter$count = 59173;
	#10 counter$count = 59174;
	#10 counter$count = 59175;
	#10 counter$count = 59176;
	#10 counter$count = 59177;
	#10 counter$count = 59178;
	#10 counter$count = 59179;
	#10 counter$count = 59180;
	#10 counter$count = 59181;
	#10 counter$count = 59182;
	#10 counter$count = 59183;
	#10 counter$count = 59184;
	#10 counter$count = 59185;
	#10 counter$count = 59186;
	#10 counter$count = 59187;
	#10 counter$count = 59188;
	#10 counter$count = 59189;
	#10 counter$count = 59190;
	#10 counter$count = 59191;
	#10 counter$count = 59192;
	#10 counter$count = 59193;
	#10 counter$count = 59194;
	#10 counter$count = 59195;
	#10 counter$count = 59196;
	#10 counter$count = 59197;
	#10 counter$count = 59198;
	#10 counter$count = 59199;
	#10 counter$count = 59200;
	#10 counter$count = 59201;
	#10 counter$count = 59202;
	#10 counter$count = 59203;
	#10 counter$count = 59204;
	#10 counter$count = 59205;
	#10 counter$count = 59206;
	#10 counter$count = 59207;
	#10 counter$count = 59208;
	#10 counter$count = 59209;
	#10 counter$count = 59210;
	#10 counter$count = 59211;
	#10 counter$count = 59212;
	#10 counter$count = 59213;
	#10 counter$count = 59214;
	#10 counter$count = 59215;
	#10 counter$count = 59216;
	#10 counter$count = 59217;
	#10 counter$count = 59218;
	#10 counter$count = 59219;
	#10 counter$count = 59220;
	#10 counter$count = 59221;
	#10 counter$count = 59222;
	#10 counter$count = 59223;
	#10 counter$count = 59224;
	#10 counter$count = 59225;
	#10 counter$count = 59226;
	#10 counter$count = 59227;
	#10 counter$count = 59228;
	#10 counter$count = 59229;
	#10 counter$count = 59230;
	#10 counter$count = 59231;
	#10 counter$count = 59232;
	#10 counter$count = 59233;
	#10 counter$count = 59234;
	#10 counter$count = 59235;
	#10 counter$count = 59236;
	#10 counter$count = 59237;
	#10 counter$count = 59238;
	#10 counter$count = 59239;
	#10 counter$count = 59240;
	#10 counter$count = 59241;
	#10 counter$count = 59242;
	#10 counter$count = 59243;
	#10 counter$count = 59244;
	#10 counter$count = 59245;
	#10 counter$count = 59246;
	#10 counter$count = 59247;
	#10 counter$count = 59248;
	#10 counter$count = 59249;
	#10 counter$count = 59250;
	#10 counter$count = 59251;
	#10 counter$count = 59252;
	#10 counter$count = 59253;
	#10 counter$count = 59254;
	#10 counter$count = 59255;
	#10 counter$count = 59256;
	#10 counter$count = 59257;
	#10 counter$count = 59258;
	#10 counter$count = 59259;
	#10 counter$count = 59260;
	#10 counter$count = 59261;
	#10 counter$count = 59262;
	#10 counter$count = 59263;
	#10 counter$count = 59264;
	#10 counter$count = 59265;
	#10 counter$count = 59266;
	#10 counter$count = 59267;
	#10 counter$count = 59268;
	#10 counter$count = 59269;
	#10 counter$count = 59270;
	#10 counter$count = 59271;
	#10 counter$count = 59272;
	#10 counter$count = 59273;
	#10 counter$count = 59274;
	#10 counter$count = 59275;
	#10 counter$count = 59276;
	#10 counter$count = 59277;
	#10 counter$count = 59278;
	#10 counter$count = 59279;
	#10 counter$count = 59280;
	#10 counter$count = 59281;
	#10 counter$count = 59282;
	#10 counter$count = 59283;
	#10 counter$count = 59284;
	#10 counter$count = 59285;
	#10 counter$count = 59286;
	#10 counter$count = 59287;
	#10 counter$count = 59288;
	#10 counter$count = 59289;
	#10 counter$count = 59290;
	#10 counter$count = 59291;
	#10 counter$count = 59292;
	#10 counter$count = 59293;
	#10 counter$count = 59294;
	#10 counter$count = 59295;
	#10 counter$count = 59296;
	#10 counter$count = 59297;
	#10 counter$count = 59298;
	#10 counter$count = 59299;
	#10 counter$count = 59300;
	#10 counter$count = 59301;
	#10 counter$count = 59302;
	#10 counter$count = 59303;
	#10 counter$count = 59304;
	#10 counter$count = 59305;
	#10 counter$count = 59306;
	#10 counter$count = 59307;
	#10 counter$count = 59308;
	#10 counter$count = 59309;
	#10 counter$count = 59310;
	#10 counter$count = 59311;
	#10 counter$count = 59312;
	#10 counter$count = 59313;
	#10 counter$count = 59314;
	#10 counter$count = 59315;
	#10 counter$count = 59316;
	#10 counter$count = 59317;
	#10 counter$count = 59318;
	#10 counter$count = 59319;
	#10 counter$count = 59320;
	#10 counter$count = 59321;
	#10 counter$count = 59322;
	#10 counter$count = 59323;
	#10 counter$count = 59324;
	#10 counter$count = 59325;
	#10 counter$count = 59326;
	#10 counter$count = 59327;
	#10 counter$count = 59328;
	#10 counter$count = 59329;
	#10 counter$count = 59330;
	#10 counter$count = 59331;
	#10 counter$count = 59332;
	#10 counter$count = 59333;
	#10 counter$count = 59334;
	#10 counter$count = 59335;
	#10 counter$count = 59336;
	#10 counter$count = 59337;
	#10 counter$count = 59338;
	#10 counter$count = 59339;
	#10 counter$count = 59340;
	#10 counter$count = 59341;
	#10 counter$count = 59342;
	#10 counter$count = 59343;
	#10 counter$count = 59344;
	#10 counter$count = 59345;
	#10 counter$count = 59346;
	#10 counter$count = 59347;
	#10 counter$count = 59348;
	#10 counter$count = 59349;
	#10 counter$count = 59350;
	#10 counter$count = 59351;
	#10 counter$count = 59352;
	#10 counter$count = 59353;
	#10 counter$count = 59354;
	#10 counter$count = 59355;
	#10 counter$count = 59356;
	#10 counter$count = 59357;
	#10 counter$count = 59358;
	#10 counter$count = 59359;
	#10 counter$count = 59360;
	#10 counter$count = 59361;
	#10 counter$count = 59362;
	#10 counter$count = 59363;
	#10 counter$count = 59364;
	#10 counter$count = 59365;
	#10 counter$count = 59366;
	#10 counter$count = 59367;
	#10 counter$count = 59368;
	#10 counter$count = 59369;
	#10 counter$count = 59370;
	#10 counter$count = 59371;
	#10 counter$count = 59372;
	#10 counter$count = 59373;
	#10 counter$count = 59374;
	#10 counter$count = 59375;
	#10 counter$count = 59376;
	#10 counter$count = 59377;
	#10 counter$count = 59378;
	#10 counter$count = 59379;
	#10 counter$count = 59380;
	#10 counter$count = 59381;
	#10 counter$count = 59382;
	#10 counter$count = 59383;
	#10 counter$count = 59384;
	#10 counter$count = 59385;
	#10 counter$count = 59386;
	#10 counter$count = 59387;
	#10 counter$count = 59388;
	#10 counter$count = 59389;
	#10 counter$count = 59390;
	#10 counter$count = 59391;
	#10 counter$count = 59392;
	#10 counter$count = 59393;
	#10 counter$count = 59394;
	#10 counter$count = 59395;
	#10 counter$count = 59396;
	#10 counter$count = 59397;
	#10 counter$count = 59398;
	#10 counter$count = 59399;
	#10 counter$count = 59400;
	#10 counter$count = 59401;
	#10 counter$count = 59402;
	#10 counter$count = 59403;
	#10 counter$count = 59404;
	#10 counter$count = 59405;
	#10 counter$count = 59406;
	#10 counter$count = 59407;
	#10 counter$count = 59408;
	#10 counter$count = 59409;
	#10 counter$count = 59410;
	#10 counter$count = 59411;
	#10 counter$count = 59412;
	#10 counter$count = 59413;
	#10 counter$count = 59414;
	#10 counter$count = 59415;
	#10 counter$count = 59416;
	#10 counter$count = 59417;
	#10 counter$count = 59418;
	#10 counter$count = 59419;
	#10 counter$count = 59420;
	#10 counter$count = 59421;
	#10 counter$count = 59422;
	#10 counter$count = 59423;
	#10 counter$count = 59424;
	#10 counter$count = 59425;
	#10 counter$count = 59426;
	#10 counter$count = 59427;
	#10 counter$count = 59428;
	#10 counter$count = 59429;
	#10 counter$count = 59430;
	#10 counter$count = 59431;
	#10 counter$count = 59432;
	#10 counter$count = 59433;
	#10 counter$count = 59434;
	#10 counter$count = 59435;
	#10 counter$count = 59436;
	#10 counter$count = 59437;
	#10 counter$count = 59438;
	#10 counter$count = 59439;
	#10 counter$count = 59440;
	#10 counter$count = 59441;
	#10 counter$count = 59442;
	#10 counter$count = 59443;
	#10 counter$count = 59444;
	#10 counter$count = 59445;
	#10 counter$count = 59446;
	#10 counter$count = 59447;
	#10 counter$count = 59448;
	#10 counter$count = 59449;
	#10 counter$count = 59450;
	#10 counter$count = 59451;
	#10 counter$count = 59452;
	#10 counter$count = 59453;
	#10 counter$count = 59454;
	#10 counter$count = 59455;
	#10 counter$count = 59456;
	#10 counter$count = 59457;
	#10 counter$count = 59458;
	#10 counter$count = 59459;
	#10 counter$count = 59460;
	#10 counter$count = 59461;
	#10 counter$count = 59462;
	#10 counter$count = 59463;
	#10 counter$count = 59464;
	#10 counter$count = 59465;
	#10 counter$count = 59466;
	#10 counter$count = 59467;
	#10 counter$count = 59468;
	#10 counter$count = 59469;
	#10 counter$count = 59470;
	#10 counter$count = 59471;
	#10 counter$count = 59472;
	#10 counter$count = 59473;
	#10 counter$count = 59474;
	#10 counter$count = 59475;
	#10 counter$count = 59476;
	#10 counter$count = 59477;
	#10 counter$count = 59478;
	#10 counter$count = 59479;
	#10 counter$count = 59480;
	#10 counter$count = 59481;
	#10 counter$count = 59482;
	#10 counter$count = 59483;
	#10 counter$count = 59484;
	#10 counter$count = 59485;
	#10 counter$count = 59486;
	#10 counter$count = 59487;
	#10 counter$count = 59488;
	#10 counter$count = 59489;
	#10 counter$count = 59490;
	#10 counter$count = 59491;
	#10 counter$count = 59492;
	#10 counter$count = 59493;
	#10 counter$count = 59494;
	#10 counter$count = 59495;
	#10 counter$count = 59496;
	#10 counter$count = 59497;
	#10 counter$count = 59498;
	#10 counter$count = 59499;
	#10 counter$count = 59500;
	#10 counter$count = 59501;
	#10 counter$count = 59502;
	#10 counter$count = 59503;
	#10 counter$count = 59504;
	#10 counter$count = 59505;
	#10 counter$count = 59506;
	#10 counter$count = 59507;
	#10 counter$count = 59508;
	#10 counter$count = 59509;
	#10 counter$count = 59510;
	#10 counter$count = 59511;
	#10 counter$count = 59512;
	#10 counter$count = 59513;
	#10 counter$count = 59514;
	#10 counter$count = 59515;
	#10 counter$count = 59516;
	#10 counter$count = 59517;
	#10 counter$count = 59518;
	#10 counter$count = 59519;
	#10 counter$count = 59520;
	#10 counter$count = 59521;
	#10 counter$count = 59522;
	#10 counter$count = 59523;
	#10 counter$count = 59524;
	#10 counter$count = 59525;
	#10 counter$count = 59526;
	#10 counter$count = 59527;
	#10 counter$count = 59528;
	#10 counter$count = 59529;
	#10 counter$count = 59530;
	#10 counter$count = 59531;
	#10 counter$count = 59532;
	#10 counter$count = 59533;
	#10 counter$count = 59534;
	#10 counter$count = 59535;
	#10 counter$count = 59536;
	#10 counter$count = 59537;
	#10 counter$count = 59538;
	#10 counter$count = 59539;
	#10 counter$count = 59540;
	#10 counter$count = 59541;
	#10 counter$count = 59542;
	#10 counter$count = 59543;
	#10 counter$count = 59544;
	#10 counter$count = 59545;
	#10 counter$count = 59546;
	#10 counter$count = 59547;
	#10 counter$count = 59548;
	#10 counter$count = 59549;
	#10 counter$count = 59550;
	#10 counter$count = 59551;
	#10 counter$count = 59552;
	#10 counter$count = 59553;
	#10 counter$count = 59554;
	#10 counter$count = 59555;
	#10 counter$count = 59556;
	#10 counter$count = 59557;
	#10 counter$count = 59558;
	#10 counter$count = 59559;
	#10 counter$count = 59560;
	#10 counter$count = 59561;
	#10 counter$count = 59562;
	#10 counter$count = 59563;
	#10 counter$count = 59564;
	#10 counter$count = 59565;
	#10 counter$count = 59566;
	#10 counter$count = 59567;
	#10 counter$count = 59568;
	#10 counter$count = 59569;
	#10 counter$count = 59570;
	#10 counter$count = 59571;
	#10 counter$count = 59572;
	#10 counter$count = 59573;
	#10 counter$count = 59574;
	#10 counter$count = 59575;
	#10 counter$count = 59576;
	#10 counter$count = 59577;
	#10 counter$count = 59578;
	#10 counter$count = 59579;
	#10 counter$count = 59580;
	#10 counter$count = 59581;
	#10 counter$count = 59582;
	#10 counter$count = 59583;
	#10 counter$count = 59584;
	#10 counter$count = 59585;
	#10 counter$count = 59586;
	#10 counter$count = 59587;
	#10 counter$count = 59588;
	#10 counter$count = 59589;
	#10 counter$count = 59590;
	#10 counter$count = 59591;
	#10 counter$count = 59592;
	#10 counter$count = 59593;
	#10 counter$count = 59594;
	#10 counter$count = 59595;
	#10 counter$count = 59596;
	#10 counter$count = 59597;
	#10 counter$count = 59598;
	#10 counter$count = 59599;
	#10 counter$count = 59600;
	#10 counter$count = 59601;
	#10 counter$count = 59602;
	#10 counter$count = 59603;
	#10 counter$count = 59604;
	#10 counter$count = 59605;
	#10 counter$count = 59606;
	#10 counter$count = 59607;
	#10 counter$count = 59608;
	#10 counter$count = 59609;
	#10 counter$count = 59610;
	#10 counter$count = 59611;
	#10 counter$count = 59612;
	#10 counter$count = 59613;
	#10 counter$count = 59614;
	#10 counter$count = 59615;
	#10 counter$count = 59616;
	#10 counter$count = 59617;
	#10 counter$count = 59618;
	#10 counter$count = 59619;
	#10 counter$count = 59620;
	#10 counter$count = 59621;
	#10 counter$count = 59622;
	#10 counter$count = 59623;
	#10 counter$count = 59624;
	#10 counter$count = 59625;
	#10 counter$count = 59626;
	#10 counter$count = 59627;
	#10 counter$count = 59628;
	#10 counter$count = 59629;
	#10 counter$count = 59630;
	#10 counter$count = 59631;
	#10 counter$count = 59632;
	#10 counter$count = 59633;
	#10 counter$count = 59634;
	#10 counter$count = 59635;
	#10 counter$count = 59636;
	#10 counter$count = 59637;
	#10 counter$count = 59638;
	#10 counter$count = 59639;
	#10 counter$count = 59640;
	#10 counter$count = 59641;
	#10 counter$count = 59642;
	#10 counter$count = 59643;
	#10 counter$count = 59644;
	#10 counter$count = 59645;
	#10 counter$count = 59646;
	#10 counter$count = 59647;
	#10 counter$count = 59648;
	#10 counter$count = 59649;
	#10 counter$count = 59650;
	#10 counter$count = 59651;
	#10 counter$count = 59652;
	#10 counter$count = 59653;
	#10 counter$count = 59654;
	#10 counter$count = 59655;
	#10 counter$count = 59656;
	#10 counter$count = 59657;
	#10 counter$count = 59658;
	#10 counter$count = 59659;
	#10 counter$count = 59660;
	#10 counter$count = 59661;
	#10 counter$count = 59662;
	#10 counter$count = 59663;
	#10 counter$count = 59664;
	#10 counter$count = 59665;
	#10 counter$count = 59666;
	#10 counter$count = 59667;
	#10 counter$count = 59668;
	#10 counter$count = 59669;
	#10 counter$count = 59670;
	#10 counter$count = 59671;
	#10 counter$count = 59672;
	#10 counter$count = 59673;
	#10 counter$count = 59674;
	#10 counter$count = 59675;
	#10 counter$count = 59676;
	#10 counter$count = 59677;
	#10 counter$count = 59678;
	#10 counter$count = 59679;
	#10 counter$count = 59680;
	#10 counter$count = 59681;
	#10 counter$count = 59682;
	#10 counter$count = 59683;
	#10 counter$count = 59684;
	#10 counter$count = 59685;
	#10 counter$count = 59686;
	#10 counter$count = 59687;
	#10 counter$count = 59688;
	#10 counter$count = 59689;
	#10 counter$count = 59690;
	#10 counter$count = 59691;
	#10 counter$count = 59692;
	#10 counter$count = 59693;
	#10 counter$count = 59694;
	#10 counter$count = 59695;
	#10 counter$count = 59696;
	#10 counter$count = 59697;
	#10 counter$count = 59698;
	#10 counter$count = 59699;
	#10 counter$count = 59700;
	#10 counter$count = 59701;
	#10 counter$count = 59702;
	#10 counter$count = 59703;
	#10 counter$count = 59704;
	#10 counter$count = 59705;
	#10 counter$count = 59706;
	#10 counter$count = 59707;
	#10 counter$count = 59708;
	#10 counter$count = 59709;
	#10 counter$count = 59710;
	#10 counter$count = 59711;
	#10 counter$count = 59712;
	#10 counter$count = 59713;
	#10 counter$count = 59714;
	#10 counter$count = 59715;
	#10 counter$count = 59716;
	#10 counter$count = 59717;
	#10 counter$count = 59718;
	#10 counter$count = 59719;
	#10 counter$count = 59720;
	#10 counter$count = 59721;
	#10 counter$count = 59722;
	#10 counter$count = 59723;
	#10 counter$count = 59724;
	#10 counter$count = 59725;
	#10 counter$count = 59726;
	#10 counter$count = 59727;
	#10 counter$count = 59728;
	#10 counter$count = 59729;
	#10 counter$count = 59730;
	#10 counter$count = 59731;
	#10 counter$count = 59732;
	#10 counter$count = 59733;
	#10 counter$count = 59734;
	#10 counter$count = 59735;
	#10 counter$count = 59736;
	#10 counter$count = 59737;
	#10 counter$count = 59738;
	#10 counter$count = 59739;
	#10 counter$count = 59740;
	#10 counter$count = 59741;
	#10 counter$count = 59742;
	#10 counter$count = 59743;
	#10 counter$count = 59744;
	#10 counter$count = 59745;
	#10 counter$count = 59746;
	#10 counter$count = 59747;
	#10 counter$count = 59748;
	#10 counter$count = 59749;
	#10 counter$count = 59750;
	#10 counter$count = 59751;
	#10 counter$count = 59752;
	#10 counter$count = 59753;
	#10 counter$count = 59754;
	#10 counter$count = 59755;
	#10 counter$count = 59756;
	#10 counter$count = 59757;
	#10 counter$count = 59758;
	#10 counter$count = 59759;
	#10 counter$count = 59760;
	#10 counter$count = 59761;
	#10 counter$count = 59762;
	#10 counter$count = 59763;
	#10 counter$count = 59764;
	#10 counter$count = 59765;
	#10 counter$count = 59766;
	#10 counter$count = 59767;
	#10 counter$count = 59768;
	#10 counter$count = 59769;
	#10 counter$count = 59770;
	#10 counter$count = 59771;
	#10 counter$count = 59772;
	#10 counter$count = 59773;
	#10 counter$count = 59774;
	#10 counter$count = 59775;
	#10 counter$count = 59776;
	#10 counter$count = 59777;
	#10 counter$count = 59778;
	#10 counter$count = 59779;
	#10 counter$count = 59780;
	#10 counter$count = 59781;
	#10 counter$count = 59782;
	#10 counter$count = 59783;
	#10 counter$count = 59784;
	#10 counter$count = 59785;
	#10 counter$count = 59786;
	#10 counter$count = 59787;
	#10 counter$count = 59788;
	#10 counter$count = 59789;
	#10 counter$count = 59790;
	#10 counter$count = 59791;
	#10 counter$count = 59792;
	#10 counter$count = 59793;
	#10 counter$count = 59794;
	#10 counter$count = 59795;
	#10 counter$count = 59796;
	#10 counter$count = 59797;
	#10 counter$count = 59798;
	#10 counter$count = 59799;
	#10 counter$count = 59800;
	#10 counter$count = 59801;
	#10 counter$count = 59802;
	#10 counter$count = 59803;
	#10 counter$count = 59804;
	#10 counter$count = 59805;
	#10 counter$count = 59806;
	#10 counter$count = 59807;
	#10 counter$count = 59808;
	#10 counter$count = 59809;
	#10 counter$count = 59810;
	#10 counter$count = 59811;
	#10 counter$count = 59812;
	#10 counter$count = 59813;
	#10 counter$count = 59814;
	#10 counter$count = 59815;
	#10 counter$count = 59816;
	#10 counter$count = 59817;
	#10 counter$count = 59818;
	#10 counter$count = 59819;
	#10 counter$count = 59820;
	#10 counter$count = 59821;
	#10 counter$count = 59822;
	#10 counter$count = 59823;
	#10 counter$count = 59824;
	#10 counter$count = 59825;
	#10 counter$count = 59826;
	#10 counter$count = 59827;
	#10 counter$count = 59828;
	#10 counter$count = 59829;
	#10 counter$count = 59830;
	#10 counter$count = 59831;
	#10 counter$count = 59832;
	#10 counter$count = 59833;
	#10 counter$count = 59834;
	#10 counter$count = 59835;
	#10 counter$count = 59836;
	#10 counter$count = 59837;
	#10 counter$count = 59838;
	#10 counter$count = 59839;
	#10 counter$count = 59840;
	#10 counter$count = 59841;
	#10 counter$count = 59842;
	#10 counter$count = 59843;
	#10 counter$count = 59844;
	#10 counter$count = 59845;
	#10 counter$count = 59846;
	#10 counter$count = 59847;
	#10 counter$count = 59848;
	#10 counter$count = 59849;
	#10 counter$count = 59850;
	#10 counter$count = 59851;
	#10 counter$count = 59852;
	#10 counter$count = 59853;
	#10 counter$count = 59854;
	#10 counter$count = 59855;
	#10 counter$count = 59856;
	#10 counter$count = 59857;
	#10 counter$count = 59858;
	#10 counter$count = 59859;
	#10 counter$count = 59860;
	#10 counter$count = 59861;
	#10 counter$count = 59862;
	#10 counter$count = 59863;
	#10 counter$count = 59864;
	#10 counter$count = 59865;
	#10 counter$count = 59866;
	#10 counter$count = 59867;
	#10 counter$count = 59868;
	#10 counter$count = 59869;
	#10 counter$count = 59870;
	#10 counter$count = 59871;
	#10 counter$count = 59872;
	#10 counter$count = 59873;
	#10 counter$count = 59874;
	#10 counter$count = 59875;
	#10 counter$count = 59876;
	#10 counter$count = 59877;
	#10 counter$count = 59878;
	#10 counter$count = 59879;
	#10 counter$count = 59880;
	#10 counter$count = 59881;
	#10 counter$count = 59882;
	#10 counter$count = 59883;
	#10 counter$count = 59884;
	#10 counter$count = 59885;
	#10 counter$count = 59886;
	#10 counter$count = 59887;
	#10 counter$count = 59888;
	#10 counter$count = 59889;
	#10 counter$count = 59890;
	#10 counter$count = 59891;
	#10 counter$count = 59892;
	#10 counter$count = 59893;
	#10 counter$count = 59894;
	#10 counter$count = 59895;
	#10 counter$count = 59896;
	#10 counter$count = 59897;
	#10 counter$count = 59898;
	#10 counter$count = 59899;
	#10 counter$count = 59900;
	#10 counter$count = 59901;
	#10 counter$count = 59902;
	#10 counter$count = 59903;
	#10 counter$count = 59904;
	#10 counter$count = 59905;
	#10 counter$count = 59906;
	#10 counter$count = 59907;
	#10 counter$count = 59908;
	#10 counter$count = 59909;
	#10 counter$count = 59910;
	#10 counter$count = 59911;
	#10 counter$count = 59912;
	#10 counter$count = 59913;
	#10 counter$count = 59914;
	#10 counter$count = 59915;
	#10 counter$count = 59916;
	#10 counter$count = 59917;
	#10 counter$count = 59918;
	#10 counter$count = 59919;
	#10 counter$count = 59920;
	#10 counter$count = 59921;
	#10 counter$count = 59922;
	#10 counter$count = 59923;
	#10 counter$count = 59924;
	#10 counter$count = 59925;
	#10 counter$count = 59926;
	#10 counter$count = 59927;
	#10 counter$count = 59928;
	#10 counter$count = 59929;
	#10 counter$count = 59930;
	#10 counter$count = 59931;
	#10 counter$count = 59932;
	#10 counter$count = 59933;
	#10 counter$count = 59934;
	#10 counter$count = 59935;
	#10 counter$count = 59936;
	#10 counter$count = 59937;
	#10 counter$count = 59938;
	#10 counter$count = 59939;
	#10 counter$count = 59940;
	#10 counter$count = 59941;
	#10 counter$count = 59942;
	#10 counter$count = 59943;
	#10 counter$count = 59944;
	#10 counter$count = 59945;
	#10 counter$count = 59946;
	#10 counter$count = 59947;
	#10 counter$count = 59948;
	#10 counter$count = 59949;
	#10 counter$count = 59950;
	#10 counter$count = 59951;
	#10 counter$count = 59952;
	#10 counter$count = 59953;
	#10 counter$count = 59954;
	#10 counter$count = 59955;
	#10 counter$count = 59956;
	#10 counter$count = 59957;
	#10 counter$count = 59958;
	#10 counter$count = 59959;
	#10 counter$count = 59960;
	#10 counter$count = 59961;
	#10 counter$count = 59962;
	#10 counter$count = 59963;
	#10 counter$count = 59964;
	#10 counter$count = 59965;
	#10 counter$count = 59966;
	#10 counter$count = 59967;
	#10 counter$count = 59968;
	#10 counter$count = 59969;
	#10 counter$count = 59970;
	#10 counter$count = 59971;
	#10 counter$count = 59972;
	#10 counter$count = 59973;
	#10 counter$count = 59974;
	#10 counter$count = 59975;
	#10 counter$count = 59976;
	#10 counter$count = 59977;
	#10 counter$count = 59978;
	#10 counter$count = 59979;
	#10 counter$count = 59980;
	#10 counter$count = 59981;
	#10 counter$count = 59982;
	#10 counter$count = 59983;
	#10 counter$count = 59984;
	#10 counter$count = 59985;
	#10 counter$count = 59986;
	#10 counter$count = 59987;
	#10 counter$count = 59988;
	#10 counter$count = 59989;
	#10 counter$count = 59990;
	#10 counter$count = 59991;
	#10 counter$count = 59992;
	#10 counter$count = 59993;
	#10 counter$count = 59994;
	#10 counter$count = 59995;
	#10 counter$count = 59996;
	#10 counter$count = 59997;
	#10 counter$count = 59998;
	#10 counter$count = 59999;
	#10 counter$count = 60000;
	#10 counter$count = 60001;
	#10 counter$count = 60002;
	#10 counter$count = 60003;
	#10 counter$count = 60004;
	#10 counter$count = 60005;
	#10 counter$count = 60006;
	#10 counter$count = 60007;
	#10 counter$count = 60008;
	#10 counter$count = 60009;
	#10 counter$count = 60010;
	#10 counter$count = 60011;
	#10 counter$count = 60012;
	#10 counter$count = 60013;
	#10 counter$count = 60014;
	#10 counter$count = 60015;
	#10 counter$count = 60016;
	#10 counter$count = 60017;
	#10 counter$count = 60018;
	#10 counter$count = 60019;
	#10 counter$count = 60020;
	#10 counter$count = 60021;
	#10 counter$count = 60022;
	#10 counter$count = 60023;
	#10 counter$count = 60024;
	#10 counter$count = 60025;
	#10 counter$count = 60026;
	#10 counter$count = 60027;
	#10 counter$count = 60028;
	#10 counter$count = 60029;
	#10 counter$count = 60030;
	#10 counter$count = 60031;
	#10 counter$count = 60032;
	#10 counter$count = 60033;
	#10 counter$count = 60034;
	#10 counter$count = 60035;
	#10 counter$count = 60036;
	#10 counter$count = 60037;
	#10 counter$count = 60038;
	#10 counter$count = 60039;
	#10 counter$count = 60040;
	#10 counter$count = 60041;
	#10 counter$count = 60042;
	#10 counter$count = 60043;
	#10 counter$count = 60044;
	#10 counter$count = 60045;
	#10 counter$count = 60046;
	#10 counter$count = 60047;
	#10 counter$count = 60048;
	#10 counter$count = 60049;
	#10 counter$count = 60050;
	#10 counter$count = 60051;
	#10 counter$count = 60052;
	#10 counter$count = 60053;
	#10 counter$count = 60054;
	#10 counter$count = 60055;
	#10 counter$count = 60056;
	#10 counter$count = 60057;
	#10 counter$count = 60058;
	#10 counter$count = 60059;
	#10 counter$count = 60060;
	#10 counter$count = 60061;
	#10 counter$count = 60062;
	#10 counter$count = 60063;
	#10 counter$count = 60064;
	#10 counter$count = 60065;
	#10 counter$count = 60066;
	#10 counter$count = 60067;
	#10 counter$count = 60068;
	#10 counter$count = 60069;
	#10 counter$count = 60070;
	#10 counter$count = 60071;
	#10 counter$count = 60072;
	#10 counter$count = 60073;
	#10 counter$count = 60074;
	#10 counter$count = 60075;
	#10 counter$count = 60076;
	#10 counter$count = 60077;
	#10 counter$count = 60078;
	#10 counter$count = 60079;
	#10 counter$count = 60080;
	#10 counter$count = 60081;
	#10 counter$count = 60082;
	#10 counter$count = 60083;
	#10 counter$count = 60084;
	#10 counter$count = 60085;
	#10 counter$count = 60086;
	#10 counter$count = 60087;
	#10 counter$count = 60088;
	#10 counter$count = 60089;
	#10 counter$count = 60090;
	#10 counter$count = 60091;
	#10 counter$count = 60092;
	#10 counter$count = 60093;
	#10 counter$count = 60094;
	#10 counter$count = 60095;
	#10 counter$count = 60096;
	#10 counter$count = 60097;
	#10 counter$count = 60098;
	#10 counter$count = 60099;
	#10 counter$count = 60100;
	#10 counter$count = 60101;
	#10 counter$count = 60102;
	#10 counter$count = 60103;
	#10 counter$count = 60104;
	#10 counter$count = 60105;
	#10 counter$count = 60106;
	#10 counter$count = 60107;
	#10 counter$count = 60108;
	#10 counter$count = 60109;
	#10 counter$count = 60110;
	#10 counter$count = 60111;
	#10 counter$count = 60112;
	#10 counter$count = 60113;
	#10 counter$count = 60114;
	#10 counter$count = 60115;
	#10 counter$count = 60116;
	#10 counter$count = 60117;
	#10 counter$count = 60118;
	#10 counter$count = 60119;
	#10 counter$count = 60120;
	#10 counter$count = 60121;
	#10 counter$count = 60122;
	#10 counter$count = 60123;
	#10 counter$count = 60124;
	#10 counter$count = 60125;
	#10 counter$count = 60126;
	#10 counter$count = 60127;
	#10 counter$count = 60128;
	#10 counter$count = 60129;
	#10 counter$count = 60130;
	#10 counter$count = 60131;
	#10 counter$count = 60132;
	#10 counter$count = 60133;
	#10 counter$count = 60134;
	#10 counter$count = 60135;
	#10 counter$count = 60136;
	#10 counter$count = 60137;
	#10 counter$count = 60138;
	#10 counter$count = 60139;
	#10 counter$count = 60140;
	#10 counter$count = 60141;
	#10 counter$count = 60142;
	#10 counter$count = 60143;
	#10 counter$count = 60144;
	#10 counter$count = 60145;
	#10 counter$count = 60146;
	#10 counter$count = 60147;
	#10 counter$count = 60148;
	#10 counter$count = 60149;
	#10 counter$count = 60150;
	#10 counter$count = 60151;
	#10 counter$count = 60152;
	#10 counter$count = 60153;
	#10 counter$count = 60154;
	#10 counter$count = 60155;
	#10 counter$count = 60156;
	#10 counter$count = 60157;
	#10 counter$count = 60158;
	#10 counter$count = 60159;
	#10 counter$count = 60160;
	#10 counter$count = 60161;
	#10 counter$count = 60162;
	#10 counter$count = 60163;
	#10 counter$count = 60164;
	#10 counter$count = 60165;
	#10 counter$count = 60166;
	#10 counter$count = 60167;
	#10 counter$count = 60168;
	#10 counter$count = 60169;
	#10 counter$count = 60170;
	#10 counter$count = 60171;
	#10 counter$count = 60172;
	#10 counter$count = 60173;
	#10 counter$count = 60174;
	#10 counter$count = 60175;
	#10 counter$count = 60176;
	#10 counter$count = 60177;
	#10 counter$count = 60178;
	#10 counter$count = 60179;
	#10 counter$count = 60180;
	#10 counter$count = 60181;
	#10 counter$count = 60182;
	#10 counter$count = 60183;
	#10 counter$count = 60184;
	#10 counter$count = 60185;
	#10 counter$count = 60186;
	#10 counter$count = 60187;
	#10 counter$count = 60188;
	#10 counter$count = 60189;
	#10 counter$count = 60190;
	#10 counter$count = 60191;
	#10 counter$count = 60192;
	#10 counter$count = 60193;
	#10 counter$count = 60194;
	#10 counter$count = 60195;
	#10 counter$count = 60196;
	#10 counter$count = 60197;
	#10 counter$count = 60198;
	#10 counter$count = 60199;
	#10 counter$count = 60200;
	#10 counter$count = 60201;
	#10 counter$count = 60202;
	#10 counter$count = 60203;
	#10 counter$count = 60204;
	#10 counter$count = 60205;
	#10 counter$count = 60206;
	#10 counter$count = 60207;
	#10 counter$count = 60208;
	#10 counter$count = 60209;
	#10 counter$count = 60210;
	#10 counter$count = 60211;
	#10 counter$count = 60212;
	#10 counter$count = 60213;
	#10 counter$count = 60214;
	#10 counter$count = 60215;
	#10 counter$count = 60216;
	#10 counter$count = 60217;
	#10 counter$count = 60218;
	#10 counter$count = 60219;
	#10 counter$count = 60220;
	#10 counter$count = 60221;
	#10 counter$count = 60222;
	#10 counter$count = 60223;
	#10 counter$count = 60224;
	#10 counter$count = 60225;
	#10 counter$count = 60226;
	#10 counter$count = 60227;
	#10 counter$count = 60228;
	#10 counter$count = 60229;
	#10 counter$count = 60230;
	#10 counter$count = 60231;
	#10 counter$count = 60232;
	#10 counter$count = 60233;
	#10 counter$count = 60234;
	#10 counter$count = 60235;
	#10 counter$count = 60236;
	#10 counter$count = 60237;
	#10 counter$count = 60238;
	#10 counter$count = 60239;
	#10 counter$count = 60240;
	#10 counter$count = 60241;
	#10 counter$count = 60242;
	#10 counter$count = 60243;
	#10 counter$count = 60244;
	#10 counter$count = 60245;
	#10 counter$count = 60246;
	#10 counter$count = 60247;
	#10 counter$count = 60248;
	#10 counter$count = 60249;
	#10 counter$count = 60250;
	#10 counter$count = 60251;
	#10 counter$count = 60252;
	#10 counter$count = 60253;
	#10 counter$count = 60254;
	#10 counter$count = 60255;
	#10 counter$count = 60256;
	#10 counter$count = 60257;
	#10 counter$count = 60258;
	#10 counter$count = 60259;
	#10 counter$count = 60260;
	#10 counter$count = 60261;
	#10 counter$count = 60262;
	#10 counter$count = 60263;
	#10 counter$count = 60264;
	#10 counter$count = 60265;
	#10 counter$count = 60266;
	#10 counter$count = 60267;
	#10 counter$count = 60268;
	#10 counter$count = 60269;
	#10 counter$count = 60270;
	#10 counter$count = 60271;
	#10 counter$count = 60272;
	#10 counter$count = 60273;
	#10 counter$count = 60274;
	#10 counter$count = 60275;
	#10 counter$count = 60276;
	#10 counter$count = 60277;
	#10 counter$count = 60278;
	#10 counter$count = 60279;
	#10 counter$count = 60280;
	#10 counter$count = 60281;
	#10 counter$count = 60282;
	#10 counter$count = 60283;
	#10 counter$count = 60284;
	#10 counter$count = 60285;
	#10 counter$count = 60286;
	#10 counter$count = 60287;
	#10 counter$count = 60288;
	#10 counter$count = 60289;
	#10 counter$count = 60290;
	#10 counter$count = 60291;
	#10 counter$count = 60292;
	#10 counter$count = 60293;
	#10 counter$count = 60294;
	#10 counter$count = 60295;
	#10 counter$count = 60296;
	#10 counter$count = 60297;
	#10 counter$count = 60298;
	#10 counter$count = 60299;
	#10 counter$count = 60300;
	#10 counter$count = 60301;
	#10 counter$count = 60302;
	#10 counter$count = 60303;
	#10 counter$count = 60304;
	#10 counter$count = 60305;
	#10 counter$count = 60306;
	#10 counter$count = 60307;
	#10 counter$count = 60308;
	#10 counter$count = 60309;
	#10 counter$count = 60310;
	#10 counter$count = 60311;
	#10 counter$count = 60312;
	#10 counter$count = 60313;
	#10 counter$count = 60314;
	#10 counter$count = 60315;
	#10 counter$count = 60316;
	#10 counter$count = 60317;
	#10 counter$count = 60318;
	#10 counter$count = 60319;
	#10 counter$count = 60320;
	#10 counter$count = 60321;
	#10 counter$count = 60322;
	#10 counter$count = 60323;
	#10 counter$count = 60324;
	#10 counter$count = 60325;
	#10 counter$count = 60326;
	#10 counter$count = 60327;
	#10 counter$count = 60328;
	#10 counter$count = 60329;
	#10 counter$count = 60330;
	#10 counter$count = 60331;
	#10 counter$count = 60332;
	#10 counter$count = 60333;
	#10 counter$count = 60334;
	#10 counter$count = 60335;
	#10 counter$count = 60336;
	#10 counter$count = 60337;
	#10 counter$count = 60338;
	#10 counter$count = 60339;
	#10 counter$count = 60340;
	#10 counter$count = 60341;
	#10 counter$count = 60342;
	#10 counter$count = 60343;
	#10 counter$count = 60344;
	#10 counter$count = 60345;
	#10 counter$count = 60346;
	#10 counter$count = 60347;
	#10 counter$count = 60348;
	#10 counter$count = 60349;
	#10 counter$count = 60350;
	#10 counter$count = 60351;
	#10 counter$count = 60352;
	#10 counter$count = 60353;
	#10 counter$count = 60354;
	#10 counter$count = 60355;
	#10 counter$count = 60356;
	#10 counter$count = 60357;
	#10 counter$count = 60358;
	#10 counter$count = 60359;
	#10 counter$count = 60360;
	#10 counter$count = 60361;
	#10 counter$count = 60362;
	#10 counter$count = 60363;
	#10 counter$count = 60364;
	#10 counter$count = 60365;
	#10 counter$count = 60366;
	#10 counter$count = 60367;
	#10 counter$count = 60368;
	#10 counter$count = 60369;
	#10 counter$count = 60370;
	#10 counter$count = 60371;
	#10 counter$count = 60372;
	#10 counter$count = 60373;
	#10 counter$count = 60374;
	#10 counter$count = 60375;
	#10 counter$count = 60376;
	#10 counter$count = 60377;
	#10 counter$count = 60378;
	#10 counter$count = 60379;
	#10 counter$count = 60380;
	#10 counter$count = 60381;
	#10 counter$count = 60382;
	#10 counter$count = 60383;
	#10 counter$count = 60384;
	#10 counter$count = 60385;
	#10 counter$count = 60386;
	#10 counter$count = 60387;
	#10 counter$count = 60388;
	#10 counter$count = 60389;
	#10 counter$count = 60390;
	#10 counter$count = 60391;
	#10 counter$count = 60392;
	#10 counter$count = 60393;
	#10 counter$count = 60394;
	#10 counter$count = 60395;
	#10 counter$count = 60396;
	#10 counter$count = 60397;
	#10 counter$count = 60398;
	#10 counter$count = 60399;
	#10 counter$count = 60400;
	#10 counter$count = 60401;
	#10 counter$count = 60402;
	#10 counter$count = 60403;
	#10 counter$count = 60404;
	#10 counter$count = 60405;
	#10 counter$count = 60406;
	#10 counter$count = 60407;
	#10 counter$count = 60408;
	#10 counter$count = 60409;
	#10 counter$count = 60410;
	#10 counter$count = 60411;
	#10 counter$count = 60412;
	#10 counter$count = 60413;
	#10 counter$count = 60414;
	#10 counter$count = 60415;
	#10 counter$count = 60416;
	#10 counter$count = 60417;
	#10 counter$count = 60418;
	#10 counter$count = 60419;
	#10 counter$count = 60420;
	#10 counter$count = 60421;
	#10 counter$count = 60422;
	#10 counter$count = 60423;
	#10 counter$count = 60424;
	#10 counter$count = 60425;
	#10 counter$count = 60426;
	#10 counter$count = 60427;
	#10 counter$count = 60428;
	#10 counter$count = 60429;
	#10 counter$count = 60430;
	#10 counter$count = 60431;
	#10 counter$count = 60432;
	#10 counter$count = 60433;
	#10 counter$count = 60434;
	#10 counter$count = 60435;
	#10 counter$count = 60436;
	#10 counter$count = 60437;
	#10 counter$count = 60438;
	#10 counter$count = 60439;
	#10 counter$count = 60440;
	#10 counter$count = 60441;
	#10 counter$count = 60442;
	#10 counter$count = 60443;
	#10 counter$count = 60444;
	#10 counter$count = 60445;
	#10 counter$count = 60446;
	#10 counter$count = 60447;
	#10 counter$count = 60448;
	#10 counter$count = 60449;
	#10 counter$count = 60450;
	#10 counter$count = 60451;
	#10 counter$count = 60452;
	#10 counter$count = 60453;
	#10 counter$count = 60454;
	#10 counter$count = 60455;
	#10 counter$count = 60456;
	#10 counter$count = 60457;
	#10 counter$count = 60458;
	#10 counter$count = 60459;
	#10 counter$count = 60460;
	#10 counter$count = 60461;
	#10 counter$count = 60462;
	#10 counter$count = 60463;
	#10 counter$count = 60464;
	#10 counter$count = 60465;
	#10 counter$count = 60466;
	#10 counter$count = 60467;
	#10 counter$count = 60468;
	#10 counter$count = 60469;
	#10 counter$count = 60470;
	#10 counter$count = 60471;
	#10 counter$count = 60472;
	#10 counter$count = 60473;
	#10 counter$count = 60474;
	#10 counter$count = 60475;
	#10 counter$count = 60476;
	#10 counter$count = 60477;
	#10 counter$count = 60478;
	#10 counter$count = 60479;
	#10 counter$count = 60480;
	#10 counter$count = 60481;
	#10 counter$count = 60482;
	#10 counter$count = 60483;
	#10 counter$count = 60484;
	#10 counter$count = 60485;
	#10 counter$count = 60486;
	#10 counter$count = 60487;
	#10 counter$count = 60488;
	#10 counter$count = 60489;
	#10 counter$count = 60490;
	#10 counter$count = 60491;
	#10 counter$count = 60492;
	#10 counter$count = 60493;
	#10 counter$count = 60494;
	#10 counter$count = 60495;
	#10 counter$count = 60496;
	#10 counter$count = 60497;
	#10 counter$count = 60498;
	#10 counter$count = 60499;
	#10 counter$count = 60500;
	#10 counter$count = 60501;
	#10 counter$count = 60502;
	#10 counter$count = 60503;
	#10 counter$count = 60504;
	#10 counter$count = 60505;
	#10 counter$count = 60506;
	#10 counter$count = 60507;
	#10 counter$count = 60508;
	#10 counter$count = 60509;
	#10 counter$count = 60510;
	#10 counter$count = 60511;
	#10 counter$count = 60512;
	#10 counter$count = 60513;
	#10 counter$count = 60514;
	#10 counter$count = 60515;
	#10 counter$count = 60516;
	#10 counter$count = 60517;
	#10 counter$count = 60518;
	#10 counter$count = 60519;
	#10 counter$count = 60520;
	#10 counter$count = 60521;
	#10 counter$count = 60522;
	#10 counter$count = 60523;
	#10 counter$count = 60524;
	#10 counter$count = 60525;
	#10 counter$count = 60526;
	#10 counter$count = 60527;
	#10 counter$count = 60528;
	#10 counter$count = 60529;
	#10 counter$count = 60530;
	#10 counter$count = 60531;
	#10 counter$count = 60532;
	#10 counter$count = 60533;
	#10 counter$count = 60534;
	#10 counter$count = 60535;
	#10 counter$count = 60536;
	#10 counter$count = 60537;
	#10 counter$count = 60538;
	#10 counter$count = 60539;
	#10 counter$count = 60540;
	#10 counter$count = 60541;
	#10 counter$count = 60542;
	#10 counter$count = 60543;
	#10 counter$count = 60544;
	#10 counter$count = 60545;
	#10 counter$count = 60546;
	#10 counter$count = 60547;
	#10 counter$count = 60548;
	#10 counter$count = 60549;
	#10 counter$count = 60550;
	#10 counter$count = 60551;
	#10 counter$count = 60552;
	#10 counter$count = 60553;
	#10 counter$count = 60554;
	#10 counter$count = 60555;
	#10 counter$count = 60556;
	#10 counter$count = 60557;
	#10 counter$count = 60558;
	#10 counter$count = 60559;
	#10 counter$count = 60560;
	#10 counter$count = 60561;
	#10 counter$count = 60562;
	#10 counter$count = 60563;
	#10 counter$count = 60564;
	#10 counter$count = 60565;
	#10 counter$count = 60566;
	#10 counter$count = 60567;
	#10 counter$count = 60568;
	#10 counter$count = 60569;
	#10 counter$count = 60570;
	#10 counter$count = 60571;
	#10 counter$count = 60572;
	#10 counter$count = 60573;
	#10 counter$count = 60574;
	#10 counter$count = 60575;
	#10 counter$count = 60576;
	#10 counter$count = 60577;
	#10 counter$count = 60578;
	#10 counter$count = 60579;
	#10 counter$count = 60580;
	#10 counter$count = 60581;
	#10 counter$count = 60582;
	#10 counter$count = 60583;
	#10 counter$count = 60584;
	#10 counter$count = 60585;
	#10 counter$count = 60586;
	#10 counter$count = 60587;
	#10 counter$count = 60588;
	#10 counter$count = 60589;
	#10 counter$count = 60590;
	#10 counter$count = 60591;
	#10 counter$count = 60592;
	#10 counter$count = 60593;
	#10 counter$count = 60594;
	#10 counter$count = 60595;
	#10 counter$count = 60596;
	#10 counter$count = 60597;
	#10 counter$count = 60598;
	#10 counter$count = 60599;
	#10 counter$count = 60600;
	#10 counter$count = 60601;
	#10 counter$count = 60602;
	#10 counter$count = 60603;
	#10 counter$count = 60604;
	#10 counter$count = 60605;
	#10 counter$count = 60606;
	#10 counter$count = 60607;
	#10 counter$count = 60608;
	#10 counter$count = 60609;
	#10 counter$count = 60610;
	#10 counter$count = 60611;
	#10 counter$count = 60612;
	#10 counter$count = 60613;
	#10 counter$count = 60614;
	#10 counter$count = 60615;
	#10 counter$count = 60616;
	#10 counter$count = 60617;
	#10 counter$count = 60618;
	#10 counter$count = 60619;
	#10 counter$count = 60620;
	#10 counter$count = 60621;
	#10 counter$count = 60622;
	#10 counter$count = 60623;
	#10 counter$count = 60624;
	#10 counter$count = 60625;
	#10 counter$count = 60626;
	#10 counter$count = 60627;
	#10 counter$count = 60628;
	#10 counter$count = 60629;
	#10 counter$count = 60630;
	#10 counter$count = 60631;
	#10 counter$count = 60632;
	#10 counter$count = 60633;
	#10 counter$count = 60634;
	#10 counter$count = 60635;
	#10 counter$count = 60636;
	#10 counter$count = 60637;
	#10 counter$count = 60638;
	#10 counter$count = 60639;
	#10 counter$count = 60640;
	#10 counter$count = 60641;
	#10 counter$count = 60642;
	#10 counter$count = 60643;
	#10 counter$count = 60644;
	#10 counter$count = 60645;
	#10 counter$count = 60646;
	#10 counter$count = 60647;
	#10 counter$count = 60648;
	#10 counter$count = 60649;
	#10 counter$count = 60650;
	#10 counter$count = 60651;
	#10 counter$count = 60652;
	#10 counter$count = 60653;
	#10 counter$count = 60654;
	#10 counter$count = 60655;
	#10 counter$count = 60656;
	#10 counter$count = 60657;
	#10 counter$count = 60658;
	#10 counter$count = 60659;
	#10 counter$count = 60660;
	#10 counter$count = 60661;
	#10 counter$count = 60662;
	#10 counter$count = 60663;
	#10 counter$count = 60664;
	#10 counter$count = 60665;
	#10 counter$count = 60666;
	#10 counter$count = 60667;
	#10 counter$count = 60668;
	#10 counter$count = 60669;
	#10 counter$count = 60670;
	#10 counter$count = 60671;
	#10 counter$count = 60672;
	#10 counter$count = 60673;
	#10 counter$count = 60674;
	#10 counter$count = 60675;
	#10 counter$count = 60676;
	#10 counter$count = 60677;
	#10 counter$count = 60678;
	#10 counter$count = 60679;
	#10 counter$count = 60680;
	#10 counter$count = 60681;
	#10 counter$count = 60682;
	#10 counter$count = 60683;
	#10 counter$count = 60684;
	#10 counter$count = 60685;
	#10 counter$count = 60686;
	#10 counter$count = 60687;
	#10 counter$count = 60688;
	#10 counter$count = 60689;
	#10 counter$count = 60690;
	#10 counter$count = 60691;
	#10 counter$count = 60692;
	#10 counter$count = 60693;
	#10 counter$count = 60694;
	#10 counter$count = 60695;
	#10 counter$count = 60696;
	#10 counter$count = 60697;
	#10 counter$count = 60698;
	#10 counter$count = 60699;
	#10 counter$count = 60700;
	#10 counter$count = 60701;
	#10 counter$count = 60702;
	#10 counter$count = 60703;
	#10 counter$count = 60704;
	#10 counter$count = 60705;
	#10 counter$count = 60706;
	#10 counter$count = 60707;
	#10 counter$count = 60708;
	#10 counter$count = 60709;
	#10 counter$count = 60710;
	#10 counter$count = 60711;
	#10 counter$count = 60712;
	#10 counter$count = 60713;
	#10 counter$count = 60714;
	#10 counter$count = 60715;
	#10 counter$count = 60716;
	#10 counter$count = 60717;
	#10 counter$count = 60718;
	#10 counter$count = 60719;
	#10 counter$count = 60720;
	#10 counter$count = 60721;
	#10 counter$count = 60722;
	#10 counter$count = 60723;
	#10 counter$count = 60724;
	#10 counter$count = 60725;
	#10 counter$count = 60726;
	#10 counter$count = 60727;
	#10 counter$count = 60728;
	#10 counter$count = 60729;
	#10 counter$count = 60730;
	#10 counter$count = 60731;
	#10 counter$count = 60732;
	#10 counter$count = 60733;
	#10 counter$count = 60734;
	#10 counter$count = 60735;
	#10 counter$count = 60736;
	#10 counter$count = 60737;
	#10 counter$count = 60738;
	#10 counter$count = 60739;
	#10 counter$count = 60740;
	#10 counter$count = 60741;
	#10 counter$count = 60742;
	#10 counter$count = 60743;
	#10 counter$count = 60744;
	#10 counter$count = 60745;
	#10 counter$count = 60746;
	#10 counter$count = 60747;
	#10 counter$count = 60748;
	#10 counter$count = 60749;
	#10 counter$count = 60750;
	#10 counter$count = 60751;
	#10 counter$count = 60752;
	#10 counter$count = 60753;
	#10 counter$count = 60754;
	#10 counter$count = 60755;
	#10 counter$count = 60756;
	#10 counter$count = 60757;
	#10 counter$count = 60758;
	#10 counter$count = 60759;
	#10 counter$count = 60760;
	#10 counter$count = 60761;
	#10 counter$count = 60762;
	#10 counter$count = 60763;
	#10 counter$count = 60764;
	#10 counter$count = 60765;
	#10 counter$count = 60766;
	#10 counter$count = 60767;
	#10 counter$count = 60768;
	#10 counter$count = 60769;
	#10 counter$count = 60770;
	#10 counter$count = 60771;
	#10 counter$count = 60772;
	#10 counter$count = 60773;
	#10 counter$count = 60774;
	#10 counter$count = 60775;
	#10 counter$count = 60776;
	#10 counter$count = 60777;
	#10 counter$count = 60778;
	#10 counter$count = 60779;
	#10 counter$count = 60780;
	#10 counter$count = 60781;
	#10 counter$count = 60782;
	#10 counter$count = 60783;
	#10 counter$count = 60784;
	#10 counter$count = 60785;
	#10 counter$count = 60786;
	#10 counter$count = 60787;
	#10 counter$count = 60788;
	#10 counter$count = 60789;
	#10 counter$count = 60790;
	#10 counter$count = 60791;
	#10 counter$count = 60792;
	#10 counter$count = 60793;
	#10 counter$count = 60794;
	#10 counter$count = 60795;
	#10 counter$count = 60796;
	#10 counter$count = 60797;
	#10 counter$count = 60798;
	#10 counter$count = 60799;
	#10 counter$count = 60800;
	#10 counter$count = 60801;
	#10 counter$count = 60802;
	#10 counter$count = 60803;
	#10 counter$count = 60804;
	#10 counter$count = 60805;
	#10 counter$count = 60806;
	#10 counter$count = 60807;
	#10 counter$count = 60808;
	#10 counter$count = 60809;
	#10 counter$count = 60810;
	#10 counter$count = 60811;
	#10 counter$count = 60812;
	#10 counter$count = 60813;
	#10 counter$count = 60814;
	#10 counter$count = 60815;
	#10 counter$count = 60816;
	#10 counter$count = 60817;
	#10 counter$count = 60818;
	#10 counter$count = 60819;
	#10 counter$count = 60820;
	#10 counter$count = 60821;
	#10 counter$count = 60822;
	#10 counter$count = 60823;
	#10 counter$count = 60824;
	#10 counter$count = 60825;
	#10 counter$count = 60826;
	#10 counter$count = 60827;
	#10 counter$count = 60828;
	#10 counter$count = 60829;
	#10 counter$count = 60830;
	#10 counter$count = 60831;
	#10 counter$count = 60832;
	#10 counter$count = 60833;
	#10 counter$count = 60834;
	#10 counter$count = 60835;
	#10 counter$count = 60836;
	#10 counter$count = 60837;
	#10 counter$count = 60838;
	#10 counter$count = 60839;
	#10 counter$count = 60840;
	#10 counter$count = 60841;
	#10 counter$count = 60842;
	#10 counter$count = 60843;
	#10 counter$count = 60844;
	#10 counter$count = 60845;
	#10 counter$count = 60846;
	#10 counter$count = 60847;
	#10 counter$count = 60848;
	#10 counter$count = 60849;
	#10 counter$count = 60850;
	#10 counter$count = 60851;
	#10 counter$count = 60852;
	#10 counter$count = 60853;
	#10 counter$count = 60854;
	#10 counter$count = 60855;
	#10 counter$count = 60856;
	#10 counter$count = 60857;
	#10 counter$count = 60858;
	#10 counter$count = 60859;
	#10 counter$count = 60860;
	#10 counter$count = 60861;
	#10 counter$count = 60862;
	#10 counter$count = 60863;
	#10 counter$count = 60864;
	#10 counter$count = 60865;
	#10 counter$count = 60866;
	#10 counter$count = 60867;
	#10 counter$count = 60868;
	#10 counter$count = 60869;
	#10 counter$count = 60870;
	#10 counter$count = 60871;
	#10 counter$count = 60872;
	#10 counter$count = 60873;
	#10 counter$count = 60874;
	#10 counter$count = 60875;
	#10 counter$count = 60876;
	#10 counter$count = 60877;
	#10 counter$count = 60878;
	#10 counter$count = 60879;
	#10 counter$count = 60880;
	#10 counter$count = 60881;
	#10 counter$count = 60882;
	#10 counter$count = 60883;
	#10 counter$count = 60884;
	#10 counter$count = 60885;
	#10 counter$count = 60886;
	#10 counter$count = 60887;
	#10 counter$count = 60888;
	#10 counter$count = 60889;
	#10 counter$count = 60890;
	#10 counter$count = 60891;
	#10 counter$count = 60892;
	#10 counter$count = 60893;
	#10 counter$count = 60894;
	#10 counter$count = 60895;
	#10 counter$count = 60896;
	#10 counter$count = 60897;
	#10 counter$count = 60898;
	#10 counter$count = 60899;
	#10 counter$count = 60900;
	#10 counter$count = 60901;
	#10 counter$count = 60902;
	#10 counter$count = 60903;
	#10 counter$count = 60904;
	#10 counter$count = 60905;
	#10 counter$count = 60906;
	#10 counter$count = 60907;
	#10 counter$count = 60908;
	#10 counter$count = 60909;
	#10 counter$count = 60910;
	#10 counter$count = 60911;
	#10 counter$count = 60912;
	#10 counter$count = 60913;
	#10 counter$count = 60914;
	#10 counter$count = 60915;
	#10 counter$count = 60916;
	#10 counter$count = 60917;
	#10 counter$count = 60918;
	#10 counter$count = 60919;
	#10 counter$count = 60920;
	#10 counter$count = 60921;
	#10 counter$count = 60922;
	#10 counter$count = 60923;
	#10 counter$count = 60924;
	#10 counter$count = 60925;
	#10 counter$count = 60926;
	#10 counter$count = 60927;
	#10 counter$count = 60928;
	#10 counter$count = 60929;
	#10 counter$count = 60930;
	#10 counter$count = 60931;
	#10 counter$count = 60932;
	#10 counter$count = 60933;
	#10 counter$count = 60934;
	#10 counter$count = 60935;
	#10 counter$count = 60936;
	#10 counter$count = 60937;
	#10 counter$count = 60938;
	#10 counter$count = 60939;
	#10 counter$count = 60940;
	#10 counter$count = 60941;
	#10 counter$count = 60942;
	#10 counter$count = 60943;
	#10 counter$count = 60944;
	#10 counter$count = 60945;
	#10 counter$count = 60946;
	#10 counter$count = 60947;
	#10 counter$count = 60948;
	#10 counter$count = 60949;
	#10 counter$count = 60950;
	#10 counter$count = 60951;
	#10 counter$count = 60952;
	#10 counter$count = 60953;
	#10 counter$count = 60954;
	#10 counter$count = 60955;
	#10 counter$count = 60956;
	#10 counter$count = 60957;
	#10 counter$count = 60958;
	#10 counter$count = 60959;
	#10 counter$count = 60960;
	#10 counter$count = 60961;
	#10 counter$count = 60962;
	#10 counter$count = 60963;
	#10 counter$count = 60964;
	#10 counter$count = 60965;
	#10 counter$count = 60966;
	#10 counter$count = 60967;
	#10 counter$count = 60968;
	#10 counter$count = 60969;
	#10 counter$count = 60970;
	#10 counter$count = 60971;
	#10 counter$count = 60972;
	#10 counter$count = 60973;
	#10 counter$count = 60974;
	#10 counter$count = 60975;
	#10 counter$count = 60976;
	#10 counter$count = 60977;
	#10 counter$count = 60978;
	#10 counter$count = 60979;
	#10 counter$count = 60980;
	#10 counter$count = 60981;
	#10 counter$count = 60982;
	#10 counter$count = 60983;
	#10 counter$count = 60984;
	#10 counter$count = 60985;
	#10 counter$count = 60986;
	#10 counter$count = 60987;
	#10 counter$count = 60988;
	#10 counter$count = 60989;
	#10 counter$count = 60990;
	#10 counter$count = 60991;
	#10 counter$count = 60992;
	#10 counter$count = 60993;
	#10 counter$count = 60994;
	#10 counter$count = 60995;
	#10 counter$count = 60996;
	#10 counter$count = 60997;
	#10 counter$count = 60998;
	#10 counter$count = 60999;
	#10 counter$count = 61000;
	#10 counter$count = 61001;
	#10 counter$count = 61002;
	#10 counter$count = 61003;
	#10 counter$count = 61004;
	#10 counter$count = 61005;
	#10 counter$count = 61006;
	#10 counter$count = 61007;
	#10 counter$count = 61008;
	#10 counter$count = 61009;
	#10 counter$count = 61010;
	#10 counter$count = 61011;
	#10 counter$count = 61012;
	#10 counter$count = 61013;
	#10 counter$count = 61014;
	#10 counter$count = 61015;
	#10 counter$count = 61016;
	#10 counter$count = 61017;
	#10 counter$count = 61018;
	#10 counter$count = 61019;
	#10 counter$count = 61020;
	#10 counter$count = 61021;
	#10 counter$count = 61022;
	#10 counter$count = 61023;
	#10 counter$count = 61024;
	#10 counter$count = 61025;
	#10 counter$count = 61026;
	#10 counter$count = 61027;
	#10 counter$count = 61028;
	#10 counter$count = 61029;
	#10 counter$count = 61030;
	#10 counter$count = 61031;
	#10 counter$count = 61032;
	#10 counter$count = 61033;
	#10 counter$count = 61034;
	#10 counter$count = 61035;
	#10 counter$count = 61036;
	#10 counter$count = 61037;
	#10 counter$count = 61038;
	#10 counter$count = 61039;
	#10 counter$count = 61040;
	#10 counter$count = 61041;
	#10 counter$count = 61042;
	#10 counter$count = 61043;
	#10 counter$count = 61044;
	#10 counter$count = 61045;
	#10 counter$count = 61046;
	#10 counter$count = 61047;
	#10 counter$count = 61048;
	#10 counter$count = 61049;
	#10 counter$count = 61050;
	#10 counter$count = 61051;
	#10 counter$count = 61052;
	#10 counter$count = 61053;
	#10 counter$count = 61054;
	#10 counter$count = 61055;
	#10 counter$count = 61056;
	#10 counter$count = 61057;
	#10 counter$count = 61058;
	#10 counter$count = 61059;
	#10 counter$count = 61060;
	#10 counter$count = 61061;
	#10 counter$count = 61062;
	#10 counter$count = 61063;
	#10 counter$count = 61064;
	#10 counter$count = 61065;
	#10 counter$count = 61066;
	#10 counter$count = 61067;
	#10 counter$count = 61068;
	#10 counter$count = 61069;
	#10 counter$count = 61070;
	#10 counter$count = 61071;
	#10 counter$count = 61072;
	#10 counter$count = 61073;
	#10 counter$count = 61074;
	#10 counter$count = 61075;
	#10 counter$count = 61076;
	#10 counter$count = 61077;
	#10 counter$count = 61078;
	#10 counter$count = 61079;
	#10 counter$count = 61080;
	#10 counter$count = 61081;
	#10 counter$count = 61082;
	#10 counter$count = 61083;
	#10 counter$count = 61084;
	#10 counter$count = 61085;
	#10 counter$count = 61086;
	#10 counter$count = 61087;
	#10 counter$count = 61088;
	#10 counter$count = 61089;
	#10 counter$count = 61090;
	#10 counter$count = 61091;
	#10 counter$count = 61092;
	#10 counter$count = 61093;
	#10 counter$count = 61094;
	#10 counter$count = 61095;
	#10 counter$count = 61096;
	#10 counter$count = 61097;
	#10 counter$count = 61098;
	#10 counter$count = 61099;
	#10 counter$count = 61100;
	#10 counter$count = 61101;
	#10 counter$count = 61102;
	#10 counter$count = 61103;
	#10 counter$count = 61104;
	#10 counter$count = 61105;
	#10 counter$count = 61106;
	#10 counter$count = 61107;
	#10 counter$count = 61108;
	#10 counter$count = 61109;
	#10 counter$count = 61110;
	#10 counter$count = 61111;
	#10 counter$count = 61112;
	#10 counter$count = 61113;
	#10 counter$count = 61114;
	#10 counter$count = 61115;
	#10 counter$count = 61116;
	#10 counter$count = 61117;
	#10 counter$count = 61118;
	#10 counter$count = 61119;
	#10 counter$count = 61120;
	#10 counter$count = 61121;
	#10 counter$count = 61122;
	#10 counter$count = 61123;
	#10 counter$count = 61124;
	#10 counter$count = 61125;
	#10 counter$count = 61126;
	#10 counter$count = 61127;
	#10 counter$count = 61128;
	#10 counter$count = 61129;
	#10 counter$count = 61130;
	#10 counter$count = 61131;
	#10 counter$count = 61132;
	#10 counter$count = 61133;
	#10 counter$count = 61134;
	#10 counter$count = 61135;
	#10 counter$count = 61136;
	#10 counter$count = 61137;
	#10 counter$count = 61138;
	#10 counter$count = 61139;
	#10 counter$count = 61140;
	#10 counter$count = 61141;
	#10 counter$count = 61142;
	#10 counter$count = 61143;
	#10 counter$count = 61144;
	#10 counter$count = 61145;
	#10 counter$count = 61146;
	#10 counter$count = 61147;
	#10 counter$count = 61148;
	#10 counter$count = 61149;
	#10 counter$count = 61150;
	#10 counter$count = 61151;
	#10 counter$count = 61152;
	#10 counter$count = 61153;
	#10 counter$count = 61154;
	#10 counter$count = 61155;
	#10 counter$count = 61156;
	#10 counter$count = 61157;
	#10 counter$count = 61158;
	#10 counter$count = 61159;
	#10 counter$count = 61160;
	#10 counter$count = 61161;
	#10 counter$count = 61162;
	#10 counter$count = 61163;
	#10 counter$count = 61164;
	#10 counter$count = 61165;
	#10 counter$count = 61166;
	#10 counter$count = 61167;
	#10 counter$count = 61168;
	#10 counter$count = 61169;
	#10 counter$count = 61170;
	#10 counter$count = 61171;
	#10 counter$count = 61172;
	#10 counter$count = 61173;
	#10 counter$count = 61174;
	#10 counter$count = 61175;
	#10 counter$count = 61176;
	#10 counter$count = 61177;
	#10 counter$count = 61178;
	#10 counter$count = 61179;
	#10 counter$count = 61180;
	#10 counter$count = 61181;
	#10 counter$count = 61182;
	#10 counter$count = 61183;
	#10 counter$count = 61184;
	#10 counter$count = 61185;
	#10 counter$count = 61186;
	#10 counter$count = 61187;
	#10 counter$count = 61188;
	#10 counter$count = 61189;
	#10 counter$count = 61190;
	#10 counter$count = 61191;
	#10 counter$count = 61192;
	#10 counter$count = 61193;
	#10 counter$count = 61194;
	#10 counter$count = 61195;
	#10 counter$count = 61196;
	#10 counter$count = 61197;
	#10 counter$count = 61198;
	#10 counter$count = 61199;
	#10 counter$count = 61200;
	#10 counter$count = 61201;
	#10 counter$count = 61202;
	#10 counter$count = 61203;
	#10 counter$count = 61204;
	#10 counter$count = 61205;
	#10 counter$count = 61206;
	#10 counter$count = 61207;
	#10 counter$count = 61208;
	#10 counter$count = 61209;
	#10 counter$count = 61210;
	#10 counter$count = 61211;
	#10 counter$count = 61212;
	#10 counter$count = 61213;
	#10 counter$count = 61214;
	#10 counter$count = 61215;
	#10 counter$count = 61216;
	#10 counter$count = 61217;
	#10 counter$count = 61218;
	#10 counter$count = 61219;
	#10 counter$count = 61220;
	#10 counter$count = 61221;
	#10 counter$count = 61222;
	#10 counter$count = 61223;
	#10 counter$count = 61224;
	#10 counter$count = 61225;
	#10 counter$count = 61226;
	#10 counter$count = 61227;
	#10 counter$count = 61228;
	#10 counter$count = 61229;
	#10 counter$count = 61230;
	#10 counter$count = 61231;
	#10 counter$count = 61232;
	#10 counter$count = 61233;
	#10 counter$count = 61234;
	#10 counter$count = 61235;
	#10 counter$count = 61236;
	#10 counter$count = 61237;
	#10 counter$count = 61238;
	#10 counter$count = 61239;
	#10 counter$count = 61240;
	#10 counter$count = 61241;
	#10 counter$count = 61242;
	#10 counter$count = 61243;
	#10 counter$count = 61244;
	#10 counter$count = 61245;
	#10 counter$count = 61246;
	#10 counter$count = 61247;
	#10 counter$count = 61248;
	#10 counter$count = 61249;
	#10 counter$count = 61250;
	#10 counter$count = 61251;
	#10 counter$count = 61252;
	#10 counter$count = 61253;
	#10 counter$count = 61254;
	#10 counter$count = 61255;
	#10 counter$count = 61256;
	#10 counter$count = 61257;
	#10 counter$count = 61258;
	#10 counter$count = 61259;
	#10 counter$count = 61260;
	#10 counter$count = 61261;
	#10 counter$count = 61262;
	#10 counter$count = 61263;
	#10 counter$count = 61264;
	#10 counter$count = 61265;
	#10 counter$count = 61266;
	#10 counter$count = 61267;
	#10 counter$count = 61268;
	#10 counter$count = 61269;
	#10 counter$count = 61270;
	#10 counter$count = 61271;
	#10 counter$count = 61272;
	#10 counter$count = 61273;
	#10 counter$count = 61274;
	#10 counter$count = 61275;
	#10 counter$count = 61276;
	#10 counter$count = 61277;
	#10 counter$count = 61278;
	#10 counter$count = 61279;
	#10 counter$count = 61280;
	#10 counter$count = 61281;
	#10 counter$count = 61282;
	#10 counter$count = 61283;
	#10 counter$count = 61284;
	#10 counter$count = 61285;
	#10 counter$count = 61286;
	#10 counter$count = 61287;
	#10 counter$count = 61288;
	#10 counter$count = 61289;
	#10 counter$count = 61290;
	#10 counter$count = 61291;
	#10 counter$count = 61292;
	#10 counter$count = 61293;
	#10 counter$count = 61294;
	#10 counter$count = 61295;
	#10 counter$count = 61296;
	#10 counter$count = 61297;
	#10 counter$count = 61298;
	#10 counter$count = 61299;
	#10 counter$count = 61300;
	#10 counter$count = 61301;
	#10 counter$count = 61302;
	#10 counter$count = 61303;
	#10 counter$count = 61304;
	#10 counter$count = 61305;
	#10 counter$count = 61306;
	#10 counter$count = 61307;
	#10 counter$count = 61308;
	#10 counter$count = 61309;
	#10 counter$count = 61310;
	#10 counter$count = 61311;
	#10 counter$count = 61312;
	#10 counter$count = 61313;
	#10 counter$count = 61314;
	#10 counter$count = 61315;
	#10 counter$count = 61316;
	#10 counter$count = 61317;
	#10 counter$count = 61318;
	#10 counter$count = 61319;
	#10 counter$count = 61320;
	#10 counter$count = 61321;
	#10 counter$count = 61322;
	#10 counter$count = 61323;
	#10 counter$count = 61324;
	#10 counter$count = 61325;
	#10 counter$count = 61326;
	#10 counter$count = 61327;
	#10 counter$count = 61328;
	#10 counter$count = 61329;
	#10 counter$count = 61330;
	#10 counter$count = 61331;
	#10 counter$count = 61332;
	#10 counter$count = 61333;
	#10 counter$count = 61334;
	#10 counter$count = 61335;
	#10 counter$count = 61336;
	#10 counter$count = 61337;
	#10 counter$count = 61338;
	#10 counter$count = 61339;
	#10 counter$count = 61340;
	#10 counter$count = 61341;
	#10 counter$count = 61342;
	#10 counter$count = 61343;
	#10 counter$count = 61344;
	#10 counter$count = 61345;
	#10 counter$count = 61346;
	#10 counter$count = 61347;
	#10 counter$count = 61348;
	#10 counter$count = 61349;
	#10 counter$count = 61350;
	#10 counter$count = 61351;
	#10 counter$count = 61352;
	#10 counter$count = 61353;
	#10 counter$count = 61354;
	#10 counter$count = 61355;
	#10 counter$count = 61356;
	#10 counter$count = 61357;
	#10 counter$count = 61358;
	#10 counter$count = 61359;
	#10 counter$count = 61360;
	#10 counter$count = 61361;
	#10 counter$count = 61362;
	#10 counter$count = 61363;
	#10 counter$count = 61364;
	#10 counter$count = 61365;
	#10 counter$count = 61366;
	#10 counter$count = 61367;
	#10 counter$count = 61368;
	#10 counter$count = 61369;
	#10 counter$count = 61370;
	#10 counter$count = 61371;
	#10 counter$count = 61372;
	#10 counter$count = 61373;
	#10 counter$count = 61374;
	#10 counter$count = 61375;
	#10 counter$count = 61376;
	#10 counter$count = 61377;
	#10 counter$count = 61378;
	#10 counter$count = 61379;
	#10 counter$count = 61380;
	#10 counter$count = 61381;
	#10 counter$count = 61382;
	#10 counter$count = 61383;
	#10 counter$count = 61384;
	#10 counter$count = 61385;
	#10 counter$count = 61386;
	#10 counter$count = 61387;
	#10 counter$count = 61388;
	#10 counter$count = 61389;
	#10 counter$count = 61390;
	#10 counter$count = 61391;
	#10 counter$count = 61392;
	#10 counter$count = 61393;
	#10 counter$count = 61394;
	#10 counter$count = 61395;
	#10 counter$count = 61396;
	#10 counter$count = 61397;
	#10 counter$count = 61398;
	#10 counter$count = 61399;
	#10 counter$count = 61400;
	#10 counter$count = 61401;
	#10 counter$count = 61402;
	#10 counter$count = 61403;
	#10 counter$count = 61404;
	#10 counter$count = 61405;
	#10 counter$count = 61406;
	#10 counter$count = 61407;
	#10 counter$count = 61408;
	#10 counter$count = 61409;
	#10 counter$count = 61410;
	#10 counter$count = 61411;
	#10 counter$count = 61412;
	#10 counter$count = 61413;
	#10 counter$count = 61414;
	#10 counter$count = 61415;
	#10 counter$count = 61416;
	#10 counter$count = 61417;
	#10 counter$count = 61418;
	#10 counter$count = 61419;
	#10 counter$count = 61420;
	#10 counter$count = 61421;
	#10 counter$count = 61422;
	#10 counter$count = 61423;
	#10 counter$count = 61424;
	#10 counter$count = 61425;
	#10 counter$count = 61426;
	#10 counter$count = 61427;
	#10 counter$count = 61428;
	#10 counter$count = 61429;
	#10 counter$count = 61430;
	#10 counter$count = 61431;
	#10 counter$count = 61432;
	#10 counter$count = 61433;
	#10 counter$count = 61434;
	#10 counter$count = 61435;
	#10 counter$count = 61436;
	#10 counter$count = 61437;
	#10 counter$count = 61438;
	#10 counter$count = 61439;
	#10 counter$count = 61440;
	#10 counter$count = 61441;
	#10 counter$count = 61442;
	#10 counter$count = 61443;
	#10 counter$count = 61444;
	#10 counter$count = 61445;
	#10 counter$count = 61446;
	#10 counter$count = 61447;
	#10 counter$count = 61448;
	#10 counter$count = 61449;
	#10 counter$count = 61450;
	#10 counter$count = 61451;
	#10 counter$count = 61452;
	#10 counter$count = 61453;
	#10 counter$count = 61454;
	#10 counter$count = 61455;
	#10 counter$count = 61456;
	#10 counter$count = 61457;
	#10 counter$count = 61458;
	#10 counter$count = 61459;
	#10 counter$count = 61460;
	#10 counter$count = 61461;
	#10 counter$count = 61462;
	#10 counter$count = 61463;
	#10 counter$count = 61464;
	#10 counter$count = 61465;
	#10 counter$count = 61466;
	#10 counter$count = 61467;
	#10 counter$count = 61468;
	#10 counter$count = 61469;
	#10 counter$count = 61470;
	#10 counter$count = 61471;
	#10 counter$count = 61472;
	#10 counter$count = 61473;
	#10 counter$count = 61474;
	#10 counter$count = 61475;
	#10 counter$count = 61476;
	#10 counter$count = 61477;
	#10 counter$count = 61478;
	#10 counter$count = 61479;
	#10 counter$count = 61480;
	#10 counter$count = 61481;
	#10 counter$count = 61482;
	#10 counter$count = 61483;
	#10 counter$count = 61484;
	#10 counter$count = 61485;
	#10 counter$count = 61486;
	#10 counter$count = 61487;
	#10 counter$count = 61488;
	#10 counter$count = 61489;
	#10 counter$count = 61490;
	#10 counter$count = 61491;
	#10 counter$count = 61492;
	#10 counter$count = 61493;
	#10 counter$count = 61494;
	#10 counter$count = 61495;
	#10 counter$count = 61496;
	#10 counter$count = 61497;
	#10 counter$count = 61498;
	#10 counter$count = 61499;
	#10 counter$count = 61500;
	#10 counter$count = 61501;
	#10 counter$count = 61502;
	#10 counter$count = 61503;
	#10 counter$count = 61504;
	#10 counter$count = 61505;
	#10 counter$count = 61506;
	#10 counter$count = 61507;
	#10 counter$count = 61508;
	#10 counter$count = 61509;
	#10 counter$count = 61510;
	#10 counter$count = 61511;
	#10 counter$count = 61512;
	#10 counter$count = 61513;
	#10 counter$count = 61514;
	#10 counter$count = 61515;
	#10 counter$count = 61516;
	#10 counter$count = 61517;
	#10 counter$count = 61518;
	#10 counter$count = 61519;
	#10 counter$count = 61520;
	#10 counter$count = 61521;
	#10 counter$count = 61522;
	#10 counter$count = 61523;
	#10 counter$count = 61524;
	#10 counter$count = 61525;
	#10 counter$count = 61526;
	#10 counter$count = 61527;
	#10 counter$count = 61528;
	#10 counter$count = 61529;
	#10 counter$count = 61530;
	#10 counter$count = 61531;
	#10 counter$count = 61532;
	#10 counter$count = 61533;
	#10 counter$count = 61534;
	#10 counter$count = 61535;
	#10 counter$count = 61536;
	#10 counter$count = 61537;
	#10 counter$count = 61538;
	#10 counter$count = 61539;
	#10 counter$count = 61540;
	#10 counter$count = 61541;
	#10 counter$count = 61542;
	#10 counter$count = 61543;
	#10 counter$count = 61544;
	#10 counter$count = 61545;
	#10 counter$count = 61546;
	#10 counter$count = 61547;
	#10 counter$count = 61548;
	#10 counter$count = 61549;
	#10 counter$count = 61550;
	#10 counter$count = 61551;
	#10 counter$count = 61552;
	#10 counter$count = 61553;
	#10 counter$count = 61554;
	#10 counter$count = 61555;
	#10 counter$count = 61556;
	#10 counter$count = 61557;
	#10 counter$count = 61558;
	#10 counter$count = 61559;
	#10 counter$count = 61560;
	#10 counter$count = 61561;
	#10 counter$count = 61562;
	#10 counter$count = 61563;
	#10 counter$count = 61564;
	#10 counter$count = 61565;
	#10 counter$count = 61566;
	#10 counter$count = 61567;
	#10 counter$count = 61568;
	#10 counter$count = 61569;
	#10 counter$count = 61570;
	#10 counter$count = 61571;
	#10 counter$count = 61572;
	#10 counter$count = 61573;
	#10 counter$count = 61574;
	#10 counter$count = 61575;
	#10 counter$count = 61576;
	#10 counter$count = 61577;
	#10 counter$count = 61578;
	#10 counter$count = 61579;
	#10 counter$count = 61580;
	#10 counter$count = 61581;
	#10 counter$count = 61582;
	#10 counter$count = 61583;
	#10 counter$count = 61584;
	#10 counter$count = 61585;
	#10 counter$count = 61586;
	#10 counter$count = 61587;
	#10 counter$count = 61588;
	#10 counter$count = 61589;
	#10 counter$count = 61590;
	#10 counter$count = 61591;
	#10 counter$count = 61592;
	#10 counter$count = 61593;
	#10 counter$count = 61594;
	#10 counter$count = 61595;
	#10 counter$count = 61596;
	#10 counter$count = 61597;
	#10 counter$count = 61598;
	#10 counter$count = 61599;
	#10 counter$count = 61600;
	#10 counter$count = 61601;
	#10 counter$count = 61602;
	#10 counter$count = 61603;
	#10 counter$count = 61604;
	#10 counter$count = 61605;
	#10 counter$count = 61606;
	#10 counter$count = 61607;
	#10 counter$count = 61608;
	#10 counter$count = 61609;
	#10 counter$count = 61610;
	#10 counter$count = 61611;
	#10 counter$count = 61612;
	#10 counter$count = 61613;
	#10 counter$count = 61614;
	#10 counter$count = 61615;
	#10 counter$count = 61616;
	#10 counter$count = 61617;
	#10 counter$count = 61618;
	#10 counter$count = 61619;
	#10 counter$count = 61620;
	#10 counter$count = 61621;
	#10 counter$count = 61622;
	#10 counter$count = 61623;
	#10 counter$count = 61624;
	#10 counter$count = 61625;
	#10 counter$count = 61626;
	#10 counter$count = 61627;
	#10 counter$count = 61628;
	#10 counter$count = 61629;
	#10 counter$count = 61630;
	#10 counter$count = 61631;
	#10 counter$count = 61632;
	#10 counter$count = 61633;
	#10 counter$count = 61634;
	#10 counter$count = 61635;
	#10 counter$count = 61636;
	#10 counter$count = 61637;
	#10 counter$count = 61638;
	#10 counter$count = 61639;
	#10 counter$count = 61640;
	#10 counter$count = 61641;
	#10 counter$count = 61642;
	#10 counter$count = 61643;
	#10 counter$count = 61644;
	#10 counter$count = 61645;
	#10 counter$count = 61646;
	#10 counter$count = 61647;
	#10 counter$count = 61648;
	#10 counter$count = 61649;
	#10 counter$count = 61650;
	#10 counter$count = 61651;
	#10 counter$count = 61652;
	#10 counter$count = 61653;
	#10 counter$count = 61654;
	#10 counter$count = 61655;
	#10 counter$count = 61656;
	#10 counter$count = 61657;
	#10 counter$count = 61658;
	#10 counter$count = 61659;
	#10 counter$count = 61660;
	#10 counter$count = 61661;
	#10 counter$count = 61662;
	#10 counter$count = 61663;
	#10 counter$count = 61664;
	#10 counter$count = 61665;
	#10 counter$count = 61666;
	#10 counter$count = 61667;
	#10 counter$count = 61668;
	#10 counter$count = 61669;
	#10 counter$count = 61670;
	#10 counter$count = 61671;
	#10 counter$count = 61672;
	#10 counter$count = 61673;
	#10 counter$count = 61674;
	#10 counter$count = 61675;
	#10 counter$count = 61676;
	#10 counter$count = 61677;
	#10 counter$count = 61678;
	#10 counter$count = 61679;
	#10 counter$count = 61680;
	#10 counter$count = 61681;
	#10 counter$count = 61682;
	#10 counter$count = 61683;
	#10 counter$count = 61684;
	#10 counter$count = 61685;
	#10 counter$count = 61686;
	#10 counter$count = 61687;
	#10 counter$count = 61688;
	#10 counter$count = 61689;
	#10 counter$count = 61690;
	#10 counter$count = 61691;
	#10 counter$count = 61692;
	#10 counter$count = 61693;
	#10 counter$count = 61694;
	#10 counter$count = 61695;
	#10 counter$count = 61696;
	#10 counter$count = 61697;
	#10 counter$count = 61698;
	#10 counter$count = 61699;
	#10 counter$count = 61700;
	#10 counter$count = 61701;
	#10 counter$count = 61702;
	#10 counter$count = 61703;
	#10 counter$count = 61704;
	#10 counter$count = 61705;
	#10 counter$count = 61706;
	#10 counter$count = 61707;
	#10 counter$count = 61708;
	#10 counter$count = 61709;
	#10 counter$count = 61710;
	#10 counter$count = 61711;
	#10 counter$count = 61712;
	#10 counter$count = 61713;
	#10 counter$count = 61714;
	#10 counter$count = 61715;
	#10 counter$count = 61716;
	#10 counter$count = 61717;
	#10 counter$count = 61718;
	#10 counter$count = 61719;
	#10 counter$count = 61720;
	#10 counter$count = 61721;
	#10 counter$count = 61722;
	#10 counter$count = 61723;
	#10 counter$count = 61724;
	#10 counter$count = 61725;
	#10 counter$count = 61726;
	#10 counter$count = 61727;
	#10 counter$count = 61728;
	#10 counter$count = 61729;
	#10 counter$count = 61730;
	#10 counter$count = 61731;
	#10 counter$count = 61732;
	#10 counter$count = 61733;
	#10 counter$count = 61734;
	#10 counter$count = 61735;
	#10 counter$count = 61736;
	#10 counter$count = 61737;
	#10 counter$count = 61738;
	#10 counter$count = 61739;
	#10 counter$count = 61740;
	#10 counter$count = 61741;
	#10 counter$count = 61742;
	#10 counter$count = 61743;
	#10 counter$count = 61744;
	#10 counter$count = 61745;
	#10 counter$count = 61746;
	#10 counter$count = 61747;
	#10 counter$count = 61748;
	#10 counter$count = 61749;
	#10 counter$count = 61750;
	#10 counter$count = 61751;
	#10 counter$count = 61752;
	#10 counter$count = 61753;
	#10 counter$count = 61754;
	#10 counter$count = 61755;
	#10 counter$count = 61756;
	#10 counter$count = 61757;
	#10 counter$count = 61758;
	#10 counter$count = 61759;
	#10 counter$count = 61760;
	#10 counter$count = 61761;
	#10 counter$count = 61762;
	#10 counter$count = 61763;
	#10 counter$count = 61764;
	#10 counter$count = 61765;
	#10 counter$count = 61766;
	#10 counter$count = 61767;
	#10 counter$count = 61768;
	#10 counter$count = 61769;
	#10 counter$count = 61770;
	#10 counter$count = 61771;
	#10 counter$count = 61772;
	#10 counter$count = 61773;
	#10 counter$count = 61774;
	#10 counter$count = 61775;
	#10 counter$count = 61776;
	#10 counter$count = 61777;
	#10 counter$count = 61778;
	#10 counter$count = 61779;
	#10 counter$count = 61780;
	#10 counter$count = 61781;
	#10 counter$count = 61782;
	#10 counter$count = 61783;
	#10 counter$count = 61784;
	#10 counter$count = 61785;
	#10 counter$count = 61786;
	#10 counter$count = 61787;
	#10 counter$count = 61788;
	#10 counter$count = 61789;
	#10 counter$count = 61790;
	#10 counter$count = 61791;
	#10 counter$count = 61792;
	#10 counter$count = 61793;
	#10 counter$count = 61794;
	#10 counter$count = 61795;
	#10 counter$count = 61796;
	#10 counter$count = 61797;
	#10 counter$count = 61798;
	#10 counter$count = 61799;
	#10 counter$count = 61800;
	#10 counter$count = 61801;
	#10 counter$count = 61802;
	#10 counter$count = 61803;
	#10 counter$count = 61804;
	#10 counter$count = 61805;
	#10 counter$count = 61806;
	#10 counter$count = 61807;
	#10 counter$count = 61808;
	#10 counter$count = 61809;
	#10 counter$count = 61810;
	#10 counter$count = 61811;
	#10 counter$count = 61812;
	#10 counter$count = 61813;
	#10 counter$count = 61814;
	#10 counter$count = 61815;
	#10 counter$count = 61816;
	#10 counter$count = 61817;
	#10 counter$count = 61818;
	#10 counter$count = 61819;
	#10 counter$count = 61820;
	#10 counter$count = 61821;
	#10 counter$count = 61822;
	#10 counter$count = 61823;
	#10 counter$count = 61824;
	#10 counter$count = 61825;
	#10 counter$count = 61826;
	#10 counter$count = 61827;
	#10 counter$count = 61828;
	#10 counter$count = 61829;
	#10 counter$count = 61830;
	#10 counter$count = 61831;
	#10 counter$count = 61832;
	#10 counter$count = 61833;
	#10 counter$count = 61834;
	#10 counter$count = 61835;
	#10 counter$count = 61836;
	#10 counter$count = 61837;
	#10 counter$count = 61838;
	#10 counter$count = 61839;
	#10 counter$count = 61840;
	#10 counter$count = 61841;
	#10 counter$count = 61842;
	#10 counter$count = 61843;
	#10 counter$count = 61844;
	#10 counter$count = 61845;
	#10 counter$count = 61846;
	#10 counter$count = 61847;
	#10 counter$count = 61848;
	#10 counter$count = 61849;
	#10 counter$count = 61850;
	#10 counter$count = 61851;
	#10 counter$count = 61852;
	#10 counter$count = 61853;
	#10 counter$count = 61854;
	#10 counter$count = 61855;
	#10 counter$count = 61856;
	#10 counter$count = 61857;
	#10 counter$count = 61858;
	#10 counter$count = 61859;
	#10 counter$count = 61860;
	#10 counter$count = 61861;
	#10 counter$count = 61862;
	#10 counter$count = 61863;
	#10 counter$count = 61864;
	#10 counter$count = 61865;
	#10 counter$count = 61866;
	#10 counter$count = 61867;
	#10 counter$count = 61868;
	#10 counter$count = 61869;
	#10 counter$count = 61870;
	#10 counter$count = 61871;
	#10 counter$count = 61872;
	#10 counter$count = 61873;
	#10 counter$count = 61874;
	#10 counter$count = 61875;
	#10 counter$count = 61876;
	#10 counter$count = 61877;
	#10 counter$count = 61878;
	#10 counter$count = 61879;
	#10 counter$count = 61880;
	#10 counter$count = 61881;
	#10 counter$count = 61882;
	#10 counter$count = 61883;
	#10 counter$count = 61884;
	#10 counter$count = 61885;
	#10 counter$count = 61886;
	#10 counter$count = 61887;
	#10 counter$count = 61888;
	#10 counter$count = 61889;
	#10 counter$count = 61890;
	#10 counter$count = 61891;
	#10 counter$count = 61892;
	#10 counter$count = 61893;
	#10 counter$count = 61894;
	#10 counter$count = 61895;
	#10 counter$count = 61896;
	#10 counter$count = 61897;
	#10 counter$count = 61898;
	#10 counter$count = 61899;
	#10 counter$count = 61900;
	#10 counter$count = 61901;
	#10 counter$count = 61902;
	#10 counter$count = 61903;
	#10 counter$count = 61904;
	#10 counter$count = 61905;
	#10 counter$count = 61906;
	#10 counter$count = 61907;
	#10 counter$count = 61908;
	#10 counter$count = 61909;
	#10 counter$count = 61910;
	#10 counter$count = 61911;
	#10 counter$count = 61912;
	#10 counter$count = 61913;
	#10 counter$count = 61914;
	#10 counter$count = 61915;
	#10 counter$count = 61916;
	#10 counter$count = 61917;
	#10 counter$count = 61918;
	#10 counter$count = 61919;
	#10 counter$count = 61920;
	#10 counter$count = 61921;
	#10 counter$count = 61922;
	#10 counter$count = 61923;
	#10 counter$count = 61924;
	#10 counter$count = 61925;
	#10 counter$count = 61926;
	#10 counter$count = 61927;
	#10 counter$count = 61928;
	#10 counter$count = 61929;
	#10 counter$count = 61930;
	#10 counter$count = 61931;
	#10 counter$count = 61932;
	#10 counter$count = 61933;
	#10 counter$count = 61934;
	#10 counter$count = 61935;
	#10 counter$count = 61936;
	#10 counter$count = 61937;
	#10 counter$count = 61938;
	#10 counter$count = 61939;
	#10 counter$count = 61940;
	#10 counter$count = 61941;
	#10 counter$count = 61942;
	#10 counter$count = 61943;
	#10 counter$count = 61944;
	#10 counter$count = 61945;
	#10 counter$count = 61946;
	#10 counter$count = 61947;
	#10 counter$count = 61948;
	#10 counter$count = 61949;
	#10 counter$count = 61950;
	#10 counter$count = 61951;
	#10 counter$count = 61952;
	#10 counter$count = 61953;
	#10 counter$count = 61954;
	#10 counter$count = 61955;
	#10 counter$count = 61956;
	#10 counter$count = 61957;
	#10 counter$count = 61958;
	#10 counter$count = 61959;
	#10 counter$count = 61960;
	#10 counter$count = 61961;
	#10 counter$count = 61962;
	#10 counter$count = 61963;
	#10 counter$count = 61964;
	#10 counter$count = 61965;
	#10 counter$count = 61966;
	#10 counter$count = 61967;
	#10 counter$count = 61968;
	#10 counter$count = 61969;
	#10 counter$count = 61970;
	#10 counter$count = 61971;
	#10 counter$count = 61972;
	#10 counter$count = 61973;
	#10 counter$count = 61974;
	#10 counter$count = 61975;
	#10 counter$count = 61976;
	#10 counter$count = 61977;
	#10 counter$count = 61978;
	#10 counter$count = 61979;
	#10 counter$count = 61980;
	#10 counter$count = 61981;
	#10 counter$count = 61982;
	#10 counter$count = 61983;
	#10 counter$count = 61984;
	#10 counter$count = 61985;
	#10 counter$count = 61986;
	#10 counter$count = 61987;
	#10 counter$count = 61988;
	#10 counter$count = 61989;
	#10 counter$count = 61990;
	#10 counter$count = 61991;
	#10 counter$count = 61992;
	#10 counter$count = 61993;
	#10 counter$count = 61994;
	#10 counter$count = 61995;
	#10 counter$count = 61996;
	#10 counter$count = 61997;
	#10 counter$count = 61998;
	#10 counter$count = 61999;
	#10 counter$count = 62000;
	#10 counter$count = 62001;
	#10 counter$count = 62002;
	#10 counter$count = 62003;
	#10 counter$count = 62004;
	#10 counter$count = 62005;
	#10 counter$count = 62006;
	#10 counter$count = 62007;
	#10 counter$count = 62008;
	#10 counter$count = 62009;
	#10 counter$count = 62010;
	#10 counter$count = 62011;
	#10 counter$count = 62012;
	#10 counter$count = 62013;
	#10 counter$count = 62014;
	#10 counter$count = 62015;
	#10 counter$count = 62016;
	#10 counter$count = 62017;
	#10 counter$count = 62018;
	#10 counter$count = 62019;
	#10 counter$count = 62020;
	#10 counter$count = 62021;
	#10 counter$count = 62022;
	#10 counter$count = 62023;
	#10 counter$count = 62024;
	#10 counter$count = 62025;
	#10 counter$count = 62026;
	#10 counter$count = 62027;
	#10 counter$count = 62028;
	#10 counter$count = 62029;
	#10 counter$count = 62030;
	#10 counter$count = 62031;
	#10 counter$count = 62032;
	#10 counter$count = 62033;
	#10 counter$count = 62034;
	#10 counter$count = 62035;
	#10 counter$count = 62036;
	#10 counter$count = 62037;
	#10 counter$count = 62038;
	#10 counter$count = 62039;
	#10 counter$count = 62040;
	#10 counter$count = 62041;
	#10 counter$count = 62042;
	#10 counter$count = 62043;
	#10 counter$count = 62044;
	#10 counter$count = 62045;
	#10 counter$count = 62046;
	#10 counter$count = 62047;
	#10 counter$count = 62048;
	#10 counter$count = 62049;
	#10 counter$count = 62050;
	#10 counter$count = 62051;
	#10 counter$count = 62052;
	#10 counter$count = 62053;
	#10 counter$count = 62054;
	#10 counter$count = 62055;
	#10 counter$count = 62056;
	#10 counter$count = 62057;
	#10 counter$count = 62058;
	#10 counter$count = 62059;
	#10 counter$count = 62060;
	#10 counter$count = 62061;
	#10 counter$count = 62062;
	#10 counter$count = 62063;
	#10 counter$count = 62064;
	#10 counter$count = 62065;
	#10 counter$count = 62066;
	#10 counter$count = 62067;
	#10 counter$count = 62068;
	#10 counter$count = 62069;
	#10 counter$count = 62070;
	#10 counter$count = 62071;
	#10 counter$count = 62072;
	#10 counter$count = 62073;
	#10 counter$count = 62074;
	#10 counter$count = 62075;
	#10 counter$count = 62076;
	#10 counter$count = 62077;
	#10 counter$count = 62078;
	#10 counter$count = 62079;
	#10 counter$count = 62080;
	#10 counter$count = 62081;
	#10 counter$count = 62082;
	#10 counter$count = 62083;
	#10 counter$count = 62084;
	#10 counter$count = 62085;
	#10 counter$count = 62086;
	#10 counter$count = 62087;
	#10 counter$count = 62088;
	#10 counter$count = 62089;
	#10 counter$count = 62090;
	#10 counter$count = 62091;
	#10 counter$count = 62092;
	#10 counter$count = 62093;
	#10 counter$count = 62094;
	#10 counter$count = 62095;
	#10 counter$count = 62096;
	#10 counter$count = 62097;
	#10 counter$count = 62098;
	#10 counter$count = 62099;
	#10 counter$count = 62100;
	#10 counter$count = 62101;
	#10 counter$count = 62102;
	#10 counter$count = 62103;
	#10 counter$count = 62104;
	#10 counter$count = 62105;
	#10 counter$count = 62106;
	#10 counter$count = 62107;
	#10 counter$count = 62108;
	#10 counter$count = 62109;
	#10 counter$count = 62110;
	#10 counter$count = 62111;
	#10 counter$count = 62112;
	#10 counter$count = 62113;
	#10 counter$count = 62114;
	#10 counter$count = 62115;
	#10 counter$count = 62116;
	#10 counter$count = 62117;
	#10 counter$count = 62118;
	#10 counter$count = 62119;
	#10 counter$count = 62120;
	#10 counter$count = 62121;
	#10 counter$count = 62122;
	#10 counter$count = 62123;
	#10 counter$count = 62124;
	#10 counter$count = 62125;
	#10 counter$count = 62126;
	#10 counter$count = 62127;
	#10 counter$count = 62128;
	#10 counter$count = 62129;
	#10 counter$count = 62130;
	#10 counter$count = 62131;
	#10 counter$count = 62132;
	#10 counter$count = 62133;
	#10 counter$count = 62134;
	#10 counter$count = 62135;
	#10 counter$count = 62136;
	#10 counter$count = 62137;
	#10 counter$count = 62138;
	#10 counter$count = 62139;
	#10 counter$count = 62140;
	#10 counter$count = 62141;
	#10 counter$count = 62142;
	#10 counter$count = 62143;
	#10 counter$count = 62144;
	#10 counter$count = 62145;
	#10 counter$count = 62146;
	#10 counter$count = 62147;
	#10 counter$count = 62148;
	#10 counter$count = 62149;
	#10 counter$count = 62150;
	#10 counter$count = 62151;
	#10 counter$count = 62152;
	#10 counter$count = 62153;
	#10 counter$count = 62154;
	#10 counter$count = 62155;
	#10 counter$count = 62156;
	#10 counter$count = 62157;
	#10 counter$count = 62158;
	#10 counter$count = 62159;
	#10 counter$count = 62160;
	#10 counter$count = 62161;
	#10 counter$count = 62162;
	#10 counter$count = 62163;
	#10 counter$count = 62164;
	#10 counter$count = 62165;
	#10 counter$count = 62166;
	#10 counter$count = 62167;
	#10 counter$count = 62168;
	#10 counter$count = 62169;
	#10 counter$count = 62170;
	#10 counter$count = 62171;
	#10 counter$count = 62172;
	#10 counter$count = 62173;
	#10 counter$count = 62174;
	#10 counter$count = 62175;
	#10 counter$count = 62176;
	#10 counter$count = 62177;
	#10 counter$count = 62178;
	#10 counter$count = 62179;
	#10 counter$count = 62180;
	#10 counter$count = 62181;
	#10 counter$count = 62182;
	#10 counter$count = 62183;
	#10 counter$count = 62184;
	#10 counter$count = 62185;
	#10 counter$count = 62186;
	#10 counter$count = 62187;
	#10 counter$count = 62188;
	#10 counter$count = 62189;
	#10 counter$count = 62190;
	#10 counter$count = 62191;
	#10 counter$count = 62192;
	#10 counter$count = 62193;
	#10 counter$count = 62194;
	#10 counter$count = 62195;
	#10 counter$count = 62196;
	#10 counter$count = 62197;
	#10 counter$count = 62198;
	#10 counter$count = 62199;
	#10 counter$count = 62200;
	#10 counter$count = 62201;
	#10 counter$count = 62202;
	#10 counter$count = 62203;
	#10 counter$count = 62204;
	#10 counter$count = 62205;
	#10 counter$count = 62206;
	#10 counter$count = 62207;
	#10 counter$count = 62208;
	#10 counter$count = 62209;
	#10 counter$count = 62210;
	#10 counter$count = 62211;
	#10 counter$count = 62212;
	#10 counter$count = 62213;
	#10 counter$count = 62214;
	#10 counter$count = 62215;
	#10 counter$count = 62216;
	#10 counter$count = 62217;
	#10 counter$count = 62218;
	#10 counter$count = 62219;
	#10 counter$count = 62220;
	#10 counter$count = 62221;
	#10 counter$count = 62222;
	#10 counter$count = 62223;
	#10 counter$count = 62224;
	#10 counter$count = 62225;
	#10 counter$count = 62226;
	#10 counter$count = 62227;
	#10 counter$count = 62228;
	#10 counter$count = 62229;
	#10 counter$count = 62230;
	#10 counter$count = 62231;
	#10 counter$count = 62232;
	#10 counter$count = 62233;
	#10 counter$count = 62234;
	#10 counter$count = 62235;
	#10 counter$count = 62236;
	#10 counter$count = 62237;
	#10 counter$count = 62238;
	#10 counter$count = 62239;
	#10 counter$count = 62240;
	#10 counter$count = 62241;
	#10 counter$count = 62242;
	#10 counter$count = 62243;
	#10 counter$count = 62244;
	#10 counter$count = 62245;
	#10 counter$count = 62246;
	#10 counter$count = 62247;
	#10 counter$count = 62248;
	#10 counter$count = 62249;
	#10 counter$count = 62250;
	#10 counter$count = 62251;
	#10 counter$count = 62252;
	#10 counter$count = 62253;
	#10 counter$count = 62254;
	#10 counter$count = 62255;
	#10 counter$count = 62256;
	#10 counter$count = 62257;
	#10 counter$count = 62258;
	#10 counter$count = 62259;
	#10 counter$count = 62260;
	#10 counter$count = 62261;
	#10 counter$count = 62262;
	#10 counter$count = 62263;
	#10 counter$count = 62264;
	#10 counter$count = 62265;
	#10 counter$count = 62266;
	#10 counter$count = 62267;
	#10 counter$count = 62268;
	#10 counter$count = 62269;
	#10 counter$count = 62270;
	#10 counter$count = 62271;
	#10 counter$count = 62272;
	#10 counter$count = 62273;
	#10 counter$count = 62274;
	#10 counter$count = 62275;
	#10 counter$count = 62276;
	#10 counter$count = 62277;
	#10 counter$count = 62278;
	#10 counter$count = 62279;
	#10 counter$count = 62280;
	#10 counter$count = 62281;
	#10 counter$count = 62282;
	#10 counter$count = 62283;
	#10 counter$count = 62284;
	#10 counter$count = 62285;
	#10 counter$count = 62286;
	#10 counter$count = 62287;
	#10 counter$count = 62288;
	#10 counter$count = 62289;
	#10 counter$count = 62290;
	#10 counter$count = 62291;
	#10 counter$count = 62292;
	#10 counter$count = 62293;
	#10 counter$count = 62294;
	#10 counter$count = 62295;
	#10 counter$count = 62296;
	#10 counter$count = 62297;
	#10 counter$count = 62298;
	#10 counter$count = 62299;
	#10 counter$count = 62300;
	#10 counter$count = 62301;
	#10 counter$count = 62302;
	#10 counter$count = 62303;
	#10 counter$count = 62304;
	#10 counter$count = 62305;
	#10 counter$count = 62306;
	#10 counter$count = 62307;
	#10 counter$count = 62308;
	#10 counter$count = 62309;
	#10 counter$count = 62310;
	#10 counter$count = 62311;
	#10 counter$count = 62312;
	#10 counter$count = 62313;
	#10 counter$count = 62314;
	#10 counter$count = 62315;
	#10 counter$count = 62316;
	#10 counter$count = 62317;
	#10 counter$count = 62318;
	#10 counter$count = 62319;
	#10 counter$count = 62320;
	#10 counter$count = 62321;
	#10 counter$count = 62322;
	#10 counter$count = 62323;
	#10 counter$count = 62324;
	#10 counter$count = 62325;
	#10 counter$count = 62326;
	#10 counter$count = 62327;
	#10 counter$count = 62328;
	#10 counter$count = 62329;
	#10 counter$count = 62330;
	#10 counter$count = 62331;
	#10 counter$count = 62332;
	#10 counter$count = 62333;
	#10 counter$count = 62334;
	#10 counter$count = 62335;
	#10 counter$count = 62336;
	#10 counter$count = 62337;
	#10 counter$count = 62338;
	#10 counter$count = 62339;
	#10 counter$count = 62340;
	#10 counter$count = 62341;
	#10 counter$count = 62342;
	#10 counter$count = 62343;
	#10 counter$count = 62344;
	#10 counter$count = 62345;
	#10 counter$count = 62346;
	#10 counter$count = 62347;
	#10 counter$count = 62348;
	#10 counter$count = 62349;
	#10 counter$count = 62350;
	#10 counter$count = 62351;
	#10 counter$count = 62352;
	#10 counter$count = 62353;
	#10 counter$count = 62354;
	#10 counter$count = 62355;
	#10 counter$count = 62356;
	#10 counter$count = 62357;
	#10 counter$count = 62358;
	#10 counter$count = 62359;
	#10 counter$count = 62360;
	#10 counter$count = 62361;
	#10 counter$count = 62362;
	#10 counter$count = 62363;
	#10 counter$count = 62364;
	#10 counter$count = 62365;
	#10 counter$count = 62366;
	#10 counter$count = 62367;
	#10 counter$count = 62368;
	#10 counter$count = 62369;
	#10 counter$count = 62370;
	#10 counter$count = 62371;
	#10 counter$count = 62372;
	#10 counter$count = 62373;
	#10 counter$count = 62374;
	#10 counter$count = 62375;
	#10 counter$count = 62376;
	#10 counter$count = 62377;
	#10 counter$count = 62378;
	#10 counter$count = 62379;
	#10 counter$count = 62380;
	#10 counter$count = 62381;
	#10 counter$count = 62382;
	#10 counter$count = 62383;
	#10 counter$count = 62384;
	#10 counter$count = 62385;
	#10 counter$count = 62386;
	#10 counter$count = 62387;
	#10 counter$count = 62388;
	#10 counter$count = 62389;
	#10 counter$count = 62390;
	#10 counter$count = 62391;
	#10 counter$count = 62392;
	#10 counter$count = 62393;
	#10 counter$count = 62394;
	#10 counter$count = 62395;
	#10 counter$count = 62396;
	#10 counter$count = 62397;
	#10 counter$count = 62398;
	#10 counter$count = 62399;
	#10 counter$count = 62400;
	#10 counter$count = 62401;
	#10 counter$count = 62402;
	#10 counter$count = 62403;
	#10 counter$count = 62404;
	#10 counter$count = 62405;
	#10 counter$count = 62406;
	#10 counter$count = 62407;
	#10 counter$count = 62408;
	#10 counter$count = 62409;
	#10 counter$count = 62410;
	#10 counter$count = 62411;
	#10 counter$count = 62412;
	#10 counter$count = 62413;
	#10 counter$count = 62414;
	#10 counter$count = 62415;
	#10 counter$count = 62416;
	#10 counter$count = 62417;
	#10 counter$count = 62418;
	#10 counter$count = 62419;
	#10 counter$count = 62420;
	#10 counter$count = 62421;
	#10 counter$count = 62422;
	#10 counter$count = 62423;
	#10 counter$count = 62424;
	#10 counter$count = 62425;
	#10 counter$count = 62426;
	#10 counter$count = 62427;
	#10 counter$count = 62428;
	#10 counter$count = 62429;
	#10 counter$count = 62430;
	#10 counter$count = 62431;
	#10 counter$count = 62432;
	#10 counter$count = 62433;
	#10 counter$count = 62434;
	#10 counter$count = 62435;
	#10 counter$count = 62436;
	#10 counter$count = 62437;
	#10 counter$count = 62438;
	#10 counter$count = 62439;
	#10 counter$count = 62440;
	#10 counter$count = 62441;
	#10 counter$count = 62442;
	#10 counter$count = 62443;
	#10 counter$count = 62444;
	#10 counter$count = 62445;
	#10 counter$count = 62446;
	#10 counter$count = 62447;
	#10 counter$count = 62448;
	#10 counter$count = 62449;
	#10 counter$count = 62450;
	#10 counter$count = 62451;
	#10 counter$count = 62452;
	#10 counter$count = 62453;
	#10 counter$count = 62454;
	#10 counter$count = 62455;
	#10 counter$count = 62456;
	#10 counter$count = 62457;
	#10 counter$count = 62458;
	#10 counter$count = 62459;
	#10 counter$count = 62460;
	#10 counter$count = 62461;
	#10 counter$count = 62462;
	#10 counter$count = 62463;
	#10 counter$count = 62464;
	#10 counter$count = 62465;
	#10 counter$count = 62466;
	#10 counter$count = 62467;
	#10 counter$count = 62468;
	#10 counter$count = 62469;
	#10 counter$count = 62470;
	#10 counter$count = 62471;
	#10 counter$count = 62472;
	#10 counter$count = 62473;
	#10 counter$count = 62474;
	#10 counter$count = 62475;
	#10 counter$count = 62476;
	#10 counter$count = 62477;
	#10 counter$count = 62478;
	#10 counter$count = 62479;
	#10 counter$count = 62480;
	#10 counter$count = 62481;
	#10 counter$count = 62482;
	#10 counter$count = 62483;
	#10 counter$count = 62484;
	#10 counter$count = 62485;
	#10 counter$count = 62486;
	#10 counter$count = 62487;
	#10 counter$count = 62488;
	#10 counter$count = 62489;
	#10 counter$count = 62490;
	#10 counter$count = 62491;
	#10 counter$count = 62492;
	#10 counter$count = 62493;
	#10 counter$count = 62494;
	#10 counter$count = 62495;
	#10 counter$count = 62496;
	#10 counter$count = 62497;
	#10 counter$count = 62498;
	#10 counter$count = 62499;
	#10 counter$count = 62500;
	#10 counter$count = 62501;
	#10 counter$count = 62502;
	#10 counter$count = 62503;
	#10 counter$count = 62504;
	#10 counter$count = 62505;
	#10 counter$count = 62506;
	#10 counter$count = 62507;
	#10 counter$count = 62508;
	#10 counter$count = 62509;
	#10 counter$count = 62510;
	#10 counter$count = 62511;
	#10 counter$count = 62512;
	#10 counter$count = 62513;
	#10 counter$count = 62514;
	#10 counter$count = 62515;
	#10 counter$count = 62516;
	#10 counter$count = 62517;
	#10 counter$count = 62518;
	#10 counter$count = 62519;
	#10 counter$count = 62520;
	#10 counter$count = 62521;
	#10 counter$count = 62522;
	#10 counter$count = 62523;
	#10 counter$count = 62524;
	#10 counter$count = 62525;
	#10 counter$count = 62526;
	#10 counter$count = 62527;
	#10 counter$count = 62528;
	#10 counter$count = 62529;
	#10 counter$count = 62530;
	#10 counter$count = 62531;
	#10 counter$count = 62532;
	#10 counter$count = 62533;
	#10 counter$count = 62534;
	#10 counter$count = 62535;
	#10 counter$count = 62536;
	#10 counter$count = 62537;
	#10 counter$count = 62538;
	#10 counter$count = 62539;
	#10 counter$count = 62540;
	#10 counter$count = 62541;
	#10 counter$count = 62542;
	#10 counter$count = 62543;
	#10 counter$count = 62544;
	#10 counter$count = 62545;
	#10 counter$count = 62546;
	#10 counter$count = 62547;
	#10 counter$count = 62548;
	#10 counter$count = 62549;
	#10 counter$count = 62550;
	#10 counter$count = 62551;
	#10 counter$count = 62552;
	#10 counter$count = 62553;
	#10 counter$count = 62554;
	#10 counter$count = 62555;
	#10 counter$count = 62556;
	#10 counter$count = 62557;
	#10 counter$count = 62558;
	#10 counter$count = 62559;
	#10 counter$count = 62560;
	#10 counter$count = 62561;
	#10 counter$count = 62562;
	#10 counter$count = 62563;
	#10 counter$count = 62564;
	#10 counter$count = 62565;
	#10 counter$count = 62566;
	#10 counter$count = 62567;
	#10 counter$count = 62568;
	#10 counter$count = 62569;
	#10 counter$count = 62570;
	#10 counter$count = 62571;
	#10 counter$count = 62572;
	#10 counter$count = 62573;
	#10 counter$count = 62574;
	#10 counter$count = 62575;
	#10 counter$count = 62576;
	#10 counter$count = 62577;
	#10 counter$count = 62578;
	#10 counter$count = 62579;
	#10 counter$count = 62580;
	#10 counter$count = 62581;
	#10 counter$count = 62582;
	#10 counter$count = 62583;
	#10 counter$count = 62584;
	#10 counter$count = 62585;
	#10 counter$count = 62586;
	#10 counter$count = 62587;
	#10 counter$count = 62588;
	#10 counter$count = 62589;
	#10 counter$count = 62590;
	#10 counter$count = 62591;
	#10 counter$count = 62592;
	#10 counter$count = 62593;
	#10 counter$count = 62594;
	#10 counter$count = 62595;
	#10 counter$count = 62596;
	#10 counter$count = 62597;
	#10 counter$count = 62598;
	#10 counter$count = 62599;
	#10 counter$count = 62600;
	#10 counter$count = 62601;
	#10 counter$count = 62602;
	#10 counter$count = 62603;
	#10 counter$count = 62604;
	#10 counter$count = 62605;
	#10 counter$count = 62606;
	#10 counter$count = 62607;
	#10 counter$count = 62608;
	#10 counter$count = 62609;
	#10 counter$count = 62610;
	#10 counter$count = 62611;
	#10 counter$count = 62612;
	#10 counter$count = 62613;
	#10 counter$count = 62614;
	#10 counter$count = 62615;
	#10 counter$count = 62616;
	#10 counter$count = 62617;
	#10 counter$count = 62618;
	#10 counter$count = 62619;
	#10 counter$count = 62620;
	#10 counter$count = 62621;
	#10 counter$count = 62622;
	#10 counter$count = 62623;
	#10 counter$count = 62624;
	#10 counter$count = 62625;
	#10 counter$count = 62626;
	#10 counter$count = 62627;
	#10 counter$count = 62628;
	#10 counter$count = 62629;
	#10 counter$count = 62630;
	#10 counter$count = 62631;
	#10 counter$count = 62632;
	#10 counter$count = 62633;
	#10 counter$count = 62634;
	#10 counter$count = 62635;
	#10 counter$count = 62636;
	#10 counter$count = 62637;
	#10 counter$count = 62638;
	#10 counter$count = 62639;
	#10 counter$count = 62640;
	#10 counter$count = 62641;
	#10 counter$count = 62642;
	#10 counter$count = 62643;
	#10 counter$count = 62644;
	#10 counter$count = 62645;
	#10 counter$count = 62646;
	#10 counter$count = 62647;
	#10 counter$count = 62648;
	#10 counter$count = 62649;
	#10 counter$count = 62650;
	#10 counter$count = 62651;
	#10 counter$count = 62652;
	#10 counter$count = 62653;
	#10 counter$count = 62654;
	#10 counter$count = 62655;
	#10 counter$count = 62656;
	#10 counter$count = 62657;
	#10 counter$count = 62658;
	#10 counter$count = 62659;
	#10 counter$count = 62660;
	#10 counter$count = 62661;
	#10 counter$count = 62662;
	#10 counter$count = 62663;
	#10 counter$count = 62664;
	#10 counter$count = 62665;
	#10 counter$count = 62666;
	#10 counter$count = 62667;
	#10 counter$count = 62668;
	#10 counter$count = 62669;
	#10 counter$count = 62670;
	#10 counter$count = 62671;
	#10 counter$count = 62672;
	#10 counter$count = 62673;
	#10 counter$count = 62674;
	#10 counter$count = 62675;
	#10 counter$count = 62676;
	#10 counter$count = 62677;
	#10 counter$count = 62678;
	#10 counter$count = 62679;
	#10 counter$count = 62680;
	#10 counter$count = 62681;
	#10 counter$count = 62682;
	#10 counter$count = 62683;
	#10 counter$count = 62684;
	#10 counter$count = 62685;
	#10 counter$count = 62686;
	#10 counter$count = 62687;
	#10 counter$count = 62688;
	#10 counter$count = 62689;
	#10 counter$count = 62690;
	#10 counter$count = 62691;
	#10 counter$count = 62692;
	#10 counter$count = 62693;
	#10 counter$count = 62694;
	#10 counter$count = 62695;
	#10 counter$count = 62696;
	#10 counter$count = 62697;
	#10 counter$count = 62698;
	#10 counter$count = 62699;
	#10 counter$count = 62700;
	#10 counter$count = 62701;
	#10 counter$count = 62702;
	#10 counter$count = 62703;
	#10 counter$count = 62704;
	#10 counter$count = 62705;
	#10 counter$count = 62706;
	#10 counter$count = 62707;
	#10 counter$count = 62708;
	#10 counter$count = 62709;
	#10 counter$count = 62710;
	#10 counter$count = 62711;
	#10 counter$count = 62712;
	#10 counter$count = 62713;
	#10 counter$count = 62714;
	#10 counter$count = 62715;
	#10 counter$count = 62716;
	#10 counter$count = 62717;
	#10 counter$count = 62718;
	#10 counter$count = 62719;
	#10 counter$count = 62720;
	#10 counter$count = 62721;
	#10 counter$count = 62722;
	#10 counter$count = 62723;
	#10 counter$count = 62724;
	#10 counter$count = 62725;
	#10 counter$count = 62726;
	#10 counter$count = 62727;
	#10 counter$count = 62728;
	#10 counter$count = 62729;
	#10 counter$count = 62730;
	#10 counter$count = 62731;
	#10 counter$count = 62732;
	#10 counter$count = 62733;
	#10 counter$count = 62734;
	#10 counter$count = 62735;
	#10 counter$count = 62736;
	#10 counter$count = 62737;
	#10 counter$count = 62738;
	#10 counter$count = 62739;
	#10 counter$count = 62740;
	#10 counter$count = 62741;
	#10 counter$count = 62742;
	#10 counter$count = 62743;
	#10 counter$count = 62744;
	#10 counter$count = 62745;
	#10 counter$count = 62746;
	#10 counter$count = 62747;
	#10 counter$count = 62748;
	#10 counter$count = 62749;
	#10 counter$count = 62750;
	#10 counter$count = 62751;
	#10 counter$count = 62752;
	#10 counter$count = 62753;
	#10 counter$count = 62754;
	#10 counter$count = 62755;
	#10 counter$count = 62756;
	#10 counter$count = 62757;
	#10 counter$count = 62758;
	#10 counter$count = 62759;
	#10 counter$count = 62760;
	#10 counter$count = 62761;
	#10 counter$count = 62762;
	#10 counter$count = 62763;
	#10 counter$count = 62764;
	#10 counter$count = 62765;
	#10 counter$count = 62766;
	#10 counter$count = 62767;
	#10 counter$count = 62768;
	#10 counter$count = 62769;
	#10 counter$count = 62770;
	#10 counter$count = 62771;
	#10 counter$count = 62772;
	#10 counter$count = 62773;
	#10 counter$count = 62774;
	#10 counter$count = 62775;
	#10 counter$count = 62776;
	#10 counter$count = 62777;
	#10 counter$count = 62778;
	#10 counter$count = 62779;
	#10 counter$count = 62780;
	#10 counter$count = 62781;
	#10 counter$count = 62782;
	#10 counter$count = 62783;
	#10 counter$count = 62784;
	#10 counter$count = 62785;
	#10 counter$count = 62786;
	#10 counter$count = 62787;
	#10 counter$count = 62788;
	#10 counter$count = 62789;
	#10 counter$count = 62790;
	#10 counter$count = 62791;
	#10 counter$count = 62792;
	#10 counter$count = 62793;
	#10 counter$count = 62794;
	#10 counter$count = 62795;
	#10 counter$count = 62796;
	#10 counter$count = 62797;
	#10 counter$count = 62798;
	#10 counter$count = 62799;
	#10 counter$count = 62800;
	#10 counter$count = 62801;
	#10 counter$count = 62802;
	#10 counter$count = 62803;
	#10 counter$count = 62804;
	#10 counter$count = 62805;
	#10 counter$count = 62806;
	#10 counter$count = 62807;
	#10 counter$count = 62808;
	#10 counter$count = 62809;
	#10 counter$count = 62810;
	#10 counter$count = 62811;
	#10 counter$count = 62812;
	#10 counter$count = 62813;
	#10 counter$count = 62814;
	#10 counter$count = 62815;
	#10 counter$count = 62816;
	#10 counter$count = 62817;
	#10 counter$count = 62818;
	#10 counter$count = 62819;
	#10 counter$count = 62820;
	#10 counter$count = 62821;
	#10 counter$count = 62822;
	#10 counter$count = 62823;
	#10 counter$count = 62824;
	#10 counter$count = 62825;
	#10 counter$count = 62826;
	#10 counter$count = 62827;
	#10 counter$count = 62828;
	#10 counter$count = 62829;
	#10 counter$count = 62830;
	#10 counter$count = 62831;
	#10 counter$count = 62832;
	#10 counter$count = 62833;
	#10 counter$count = 62834;
	#10 counter$count = 62835;
	#10 counter$count = 62836;
	#10 counter$count = 62837;
	#10 counter$count = 62838;
	#10 counter$count = 62839;
	#10 counter$count = 62840;
	#10 counter$count = 62841;
	#10 counter$count = 62842;
	#10 counter$count = 62843;
	#10 counter$count = 62844;
	#10 counter$count = 62845;
	#10 counter$count = 62846;
	#10 counter$count = 62847;
	#10 counter$count = 62848;
	#10 counter$count = 62849;
	#10 counter$count = 62850;
	#10 counter$count = 62851;
	#10 counter$count = 62852;
	#10 counter$count = 62853;
	#10 counter$count = 62854;
	#10 counter$count = 62855;
	#10 counter$count = 62856;
	#10 counter$count = 62857;
	#10 counter$count = 62858;
	#10 counter$count = 62859;
	#10 counter$count = 62860;
	#10 counter$count = 62861;
	#10 counter$count = 62862;
	#10 counter$count = 62863;
	#10 counter$count = 62864;
	#10 counter$count = 62865;
	#10 counter$count = 62866;
	#10 counter$count = 62867;
	#10 counter$count = 62868;
	#10 counter$count = 62869;
	#10 counter$count = 62870;
	#10 counter$count = 62871;
	#10 counter$count = 62872;
	#10 counter$count = 62873;
	#10 counter$count = 62874;
	#10 counter$count = 62875;
	#10 counter$count = 62876;
	#10 counter$count = 62877;
	#10 counter$count = 62878;
	#10 counter$count = 62879;
	#10 counter$count = 62880;
	#10 counter$count = 62881;
	#10 counter$count = 62882;
	#10 counter$count = 62883;
	#10 counter$count = 62884;
	#10 counter$count = 62885;
	#10 counter$count = 62886;
	#10 counter$count = 62887;
	#10 counter$count = 62888;
	#10 counter$count = 62889;
	#10 counter$count = 62890;
	#10 counter$count = 62891;
	#10 counter$count = 62892;
	#10 counter$count = 62893;
	#10 counter$count = 62894;
	#10 counter$count = 62895;
	#10 counter$count = 62896;
	#10 counter$count = 62897;
	#10 counter$count = 62898;
	#10 counter$count = 62899;
	#10 counter$count = 62900;
	#10 counter$count = 62901;
	#10 counter$count = 62902;
	#10 counter$count = 62903;
	#10 counter$count = 62904;
	#10 counter$count = 62905;
	#10 counter$count = 62906;
	#10 counter$count = 62907;
	#10 counter$count = 62908;
	#10 counter$count = 62909;
	#10 counter$count = 62910;
	#10 counter$count = 62911;
	#10 counter$count = 62912;
	#10 counter$count = 62913;
	#10 counter$count = 62914;
	#10 counter$count = 62915;
	#10 counter$count = 62916;
	#10 counter$count = 62917;
	#10 counter$count = 62918;
	#10 counter$count = 62919;
	#10 counter$count = 62920;
	#10 counter$count = 62921;
	#10 counter$count = 62922;
	#10 counter$count = 62923;
	#10 counter$count = 62924;
	#10 counter$count = 62925;
	#10 counter$count = 62926;
	#10 counter$count = 62927;
	#10 counter$count = 62928;
	#10 counter$count = 62929;
	#10 counter$count = 62930;
	#10 counter$count = 62931;
	#10 counter$count = 62932;
	#10 counter$count = 62933;
	#10 counter$count = 62934;
	#10 counter$count = 62935;
	#10 counter$count = 62936;
	#10 counter$count = 62937;
	#10 counter$count = 62938;
	#10 counter$count = 62939;
	#10 counter$count = 62940;
	#10 counter$count = 62941;
	#10 counter$count = 62942;
	#10 counter$count = 62943;
	#10 counter$count = 62944;
	#10 counter$count = 62945;
	#10 counter$count = 62946;
	#10 counter$count = 62947;
	#10 counter$count = 62948;
	#10 counter$count = 62949;
	#10 counter$count = 62950;
	#10 counter$count = 62951;
	#10 counter$count = 62952;
	#10 counter$count = 62953;
	#10 counter$count = 62954;
	#10 counter$count = 62955;
	#10 counter$count = 62956;
	#10 counter$count = 62957;
	#10 counter$count = 62958;
	#10 counter$count = 62959;
	#10 counter$count = 62960;
	#10 counter$count = 62961;
	#10 counter$count = 62962;
	#10 counter$count = 62963;
	#10 counter$count = 62964;
	#10 counter$count = 62965;
	#10 counter$count = 62966;
	#10 counter$count = 62967;
	#10 counter$count = 62968;
	#10 counter$count = 62969;
	#10 counter$count = 62970;
	#10 counter$count = 62971;
	#10 counter$count = 62972;
	#10 counter$count = 62973;
	#10 counter$count = 62974;
	#10 counter$count = 62975;
	#10 counter$count = 62976;
	#10 counter$count = 62977;
	#10 counter$count = 62978;
	#10 counter$count = 62979;
	#10 counter$count = 62980;
	#10 counter$count = 62981;
	#10 counter$count = 62982;
	#10 counter$count = 62983;
	#10 counter$count = 62984;
	#10 counter$count = 62985;
	#10 counter$count = 62986;
	#10 counter$count = 62987;
	#10 counter$count = 62988;
	#10 counter$count = 62989;
	#10 counter$count = 62990;
	#10 counter$count = 62991;
	#10 counter$count = 62992;
	#10 counter$count = 62993;
	#10 counter$count = 62994;
	#10 counter$count = 62995;
	#10 counter$count = 62996;
	#10 counter$count = 62997;
	#10 counter$count = 62998;
	#10 counter$count = 62999;
	#10 counter$count = 63000;
	#10 counter$count = 63001;
	#10 counter$count = 63002;
	#10 counter$count = 63003;
	#10 counter$count = 63004;
	#10 counter$count = 63005;
	#10 counter$count = 63006;
	#10 counter$count = 63007;
	#10 counter$count = 63008;
	#10 counter$count = 63009;
	#10 counter$count = 63010;
	#10 counter$count = 63011;
	#10 counter$count = 63012;
	#10 counter$count = 63013;
	#10 counter$count = 63014;
	#10 counter$count = 63015;
	#10 counter$count = 63016;
	#10 counter$count = 63017;
	#10 counter$count = 63018;
	#10 counter$count = 63019;
	#10 counter$count = 63020;
	#10 counter$count = 63021;
	#10 counter$count = 63022;
	#10 counter$count = 63023;
	#10 counter$count = 63024;
	#10 counter$count = 63025;
	#10 counter$count = 63026;
	#10 counter$count = 63027;
	#10 counter$count = 63028;
	#10 counter$count = 63029;
	#10 counter$count = 63030;
	#10 counter$count = 63031;
	#10 counter$count = 63032;
	#10 counter$count = 63033;
	#10 counter$count = 63034;
	#10 counter$count = 63035;
	#10 counter$count = 63036;
	#10 counter$count = 63037;
	#10 counter$count = 63038;
	#10 counter$count = 63039;
	#10 counter$count = 63040;
	#10 counter$count = 63041;
	#10 counter$count = 63042;
	#10 counter$count = 63043;
	#10 counter$count = 63044;
	#10 counter$count = 63045;
	#10 counter$count = 63046;
	#10 counter$count = 63047;
	#10 counter$count = 63048;
	#10 counter$count = 63049;
	#10 counter$count = 63050;
	#10 counter$count = 63051;
	#10 counter$count = 63052;
	#10 counter$count = 63053;
	#10 counter$count = 63054;
	#10 counter$count = 63055;
	#10 counter$count = 63056;
	#10 counter$count = 63057;
	#10 counter$count = 63058;
	#10 counter$count = 63059;
	#10 counter$count = 63060;
	#10 counter$count = 63061;
	#10 counter$count = 63062;
	#10 counter$count = 63063;
	#10 counter$count = 63064;
	#10 counter$count = 63065;
	#10 counter$count = 63066;
	#10 counter$count = 63067;
	#10 counter$count = 63068;
	#10 counter$count = 63069;
	#10 counter$count = 63070;
	#10 counter$count = 63071;
	#10 counter$count = 63072;
	#10 counter$count = 63073;
	#10 counter$count = 63074;
	#10 counter$count = 63075;
	#10 counter$count = 63076;
	#10 counter$count = 63077;
	#10 counter$count = 63078;
	#10 counter$count = 63079;
	#10 counter$count = 63080;
	#10 counter$count = 63081;
	#10 counter$count = 63082;
	#10 counter$count = 63083;
	#10 counter$count = 63084;
	#10 counter$count = 63085;
	#10 counter$count = 63086;
	#10 counter$count = 63087;
	#10 counter$count = 63088;
	#10 counter$count = 63089;
	#10 counter$count = 63090;
	#10 counter$count = 63091;
	#10 counter$count = 63092;
	#10 counter$count = 63093;
	#10 counter$count = 63094;
	#10 counter$count = 63095;
	#10 counter$count = 63096;
	#10 counter$count = 63097;
	#10 counter$count = 63098;
	#10 counter$count = 63099;
	#10 counter$count = 63100;
	#10 counter$count = 63101;
	#10 counter$count = 63102;
	#10 counter$count = 63103;
	#10 counter$count = 63104;
	#10 counter$count = 63105;
	#10 counter$count = 63106;
	#10 counter$count = 63107;
	#10 counter$count = 63108;
	#10 counter$count = 63109;
	#10 counter$count = 63110;
	#10 counter$count = 63111;
	#10 counter$count = 63112;
	#10 counter$count = 63113;
	#10 counter$count = 63114;
	#10 counter$count = 63115;
	#10 counter$count = 63116;
	#10 counter$count = 63117;
	#10 counter$count = 63118;
	#10 counter$count = 63119;
	#10 counter$count = 63120;
	#10 counter$count = 63121;
	#10 counter$count = 63122;
	#10 counter$count = 63123;
	#10 counter$count = 63124;
	#10 counter$count = 63125;
	#10 counter$count = 63126;
	#10 counter$count = 63127;
	#10 counter$count = 63128;
	#10 counter$count = 63129;
	#10 counter$count = 63130;
	#10 counter$count = 63131;
	#10 counter$count = 63132;
	#10 counter$count = 63133;
	#10 counter$count = 63134;
	#10 counter$count = 63135;
	#10 counter$count = 63136;
	#10 counter$count = 63137;
	#10 counter$count = 63138;
	#10 counter$count = 63139;
	#10 counter$count = 63140;
	#10 counter$count = 63141;
	#10 counter$count = 63142;
	#10 counter$count = 63143;
	#10 counter$count = 63144;
	#10 counter$count = 63145;
	#10 counter$count = 63146;
	#10 counter$count = 63147;
	#10 counter$count = 63148;
	#10 counter$count = 63149;
	#10 counter$count = 63150;
	#10 counter$count = 63151;
	#10 counter$count = 63152;
	#10 counter$count = 63153;
	#10 counter$count = 63154;
	#10 counter$count = 63155;
	#10 counter$count = 63156;
	#10 counter$count = 63157;
	#10 counter$count = 63158;
	#10 counter$count = 63159;
	#10 counter$count = 63160;
	#10 counter$count = 63161;
	#10 counter$count = 63162;
	#10 counter$count = 63163;
	#10 counter$count = 63164;
	#10 counter$count = 63165;
	#10 counter$count = 63166;
	#10 counter$count = 63167;
	#10 counter$count = 63168;
	#10 counter$count = 63169;
	#10 counter$count = 63170;
	#10 counter$count = 63171;
	#10 counter$count = 63172;
	#10 counter$count = 63173;
	#10 counter$count = 63174;
	#10 counter$count = 63175;
	#10 counter$count = 63176;
	#10 counter$count = 63177;
	#10 counter$count = 63178;
	#10 counter$count = 63179;
	#10 counter$count = 63180;
	#10 counter$count = 63181;
	#10 counter$count = 63182;
	#10 counter$count = 63183;
	#10 counter$count = 63184;
	#10 counter$count = 63185;
	#10 counter$count = 63186;
	#10 counter$count = 63187;
	#10 counter$count = 63188;
	#10 counter$count = 63189;
	#10 counter$count = 63190;
	#10 counter$count = 63191;
	#10 counter$count = 63192;
	#10 counter$count = 63193;
	#10 counter$count = 63194;
	#10 counter$count = 63195;
	#10 counter$count = 63196;
	#10 counter$count = 63197;
	#10 counter$count = 63198;
	#10 counter$count = 63199;
	#10 counter$count = 63200;
	#10 counter$count = 63201;
	#10 counter$count = 63202;
	#10 counter$count = 63203;
	#10 counter$count = 63204;
	#10 counter$count = 63205;
	#10 counter$count = 63206;
	#10 counter$count = 63207;
	#10 counter$count = 63208;
	#10 counter$count = 63209;
	#10 counter$count = 63210;
	#10 counter$count = 63211;
	#10 counter$count = 63212;
	#10 counter$count = 63213;
	#10 counter$count = 63214;
	#10 counter$count = 63215;
	#10 counter$count = 63216;
	#10 counter$count = 63217;
	#10 counter$count = 63218;
	#10 counter$count = 63219;
	#10 counter$count = 63220;
	#10 counter$count = 63221;
	#10 counter$count = 63222;
	#10 counter$count = 63223;
	#10 counter$count = 63224;
	#10 counter$count = 63225;
	#10 counter$count = 63226;
	#10 counter$count = 63227;
	#10 counter$count = 63228;
	#10 counter$count = 63229;
	#10 counter$count = 63230;
	#10 counter$count = 63231;
	#10 counter$count = 63232;
	#10 counter$count = 63233;
	#10 counter$count = 63234;
	#10 counter$count = 63235;
	#10 counter$count = 63236;
	#10 counter$count = 63237;
	#10 counter$count = 63238;
	#10 counter$count = 63239;
	#10 counter$count = 63240;
	#10 counter$count = 63241;
	#10 counter$count = 63242;
	#10 counter$count = 63243;
	#10 counter$count = 63244;
	#10 counter$count = 63245;
	#10 counter$count = 63246;
	#10 counter$count = 63247;
	#10 counter$count = 63248;
	#10 counter$count = 63249;
	#10 counter$count = 63250;
	#10 counter$count = 63251;
	#10 counter$count = 63252;
	#10 counter$count = 63253;
	#10 counter$count = 63254;
	#10 counter$count = 63255;
	#10 counter$count = 63256;
	#10 counter$count = 63257;
	#10 counter$count = 63258;
	#10 counter$count = 63259;
	#10 counter$count = 63260;
	#10 counter$count = 63261;
	#10 counter$count = 63262;
	#10 counter$count = 63263;
	#10 counter$count = 63264;
	#10 counter$count = 63265;
	#10 counter$count = 63266;
	#10 counter$count = 63267;
	#10 counter$count = 63268;
	#10 counter$count = 63269;
	#10 counter$count = 63270;
	#10 counter$count = 63271;
	#10 counter$count = 63272;
	#10 counter$count = 63273;
	#10 counter$count = 63274;
	#10 counter$count = 63275;
	#10 counter$count = 63276;
	#10 counter$count = 63277;
	#10 counter$count = 63278;
	#10 counter$count = 63279;
	#10 counter$count = 63280;
	#10 counter$count = 63281;
	#10 counter$count = 63282;
	#10 counter$count = 63283;
	#10 counter$count = 63284;
	#10 counter$count = 63285;
	#10 counter$count = 63286;
	#10 counter$count = 63287;
	#10 counter$count = 63288;
	#10 counter$count = 63289;
	#10 counter$count = 63290;
	#10 counter$count = 63291;
	#10 counter$count = 63292;
	#10 counter$count = 63293;
	#10 counter$count = 63294;
	#10 counter$count = 63295;
	#10 counter$count = 63296;
	#10 counter$count = 63297;
	#10 counter$count = 63298;
	#10 counter$count = 63299;
	#10 counter$count = 63300;
	#10 counter$count = 63301;
	#10 counter$count = 63302;
	#10 counter$count = 63303;
	#10 counter$count = 63304;
	#10 counter$count = 63305;
	#10 counter$count = 63306;
	#10 counter$count = 63307;
	#10 counter$count = 63308;
	#10 counter$count = 63309;
	#10 counter$count = 63310;
	#10 counter$count = 63311;
	#10 counter$count = 63312;
	#10 counter$count = 63313;
	#10 counter$count = 63314;
	#10 counter$count = 63315;
	#10 counter$count = 63316;
	#10 counter$count = 63317;
	#10 counter$count = 63318;
	#10 counter$count = 63319;
	#10 counter$count = 63320;
	#10 counter$count = 63321;
	#10 counter$count = 63322;
	#10 counter$count = 63323;
	#10 counter$count = 63324;
	#10 counter$count = 63325;
	#10 counter$count = 63326;
	#10 counter$count = 63327;
	#10 counter$count = 63328;
	#10 counter$count = 63329;
	#10 counter$count = 63330;
	#10 counter$count = 63331;
	#10 counter$count = 63332;
	#10 counter$count = 63333;
	#10 counter$count = 63334;
	#10 counter$count = 63335;
	#10 counter$count = 63336;
	#10 counter$count = 63337;
	#10 counter$count = 63338;
	#10 counter$count = 63339;
	#10 counter$count = 63340;
	#10 counter$count = 63341;
	#10 counter$count = 63342;
	#10 counter$count = 63343;
	#10 counter$count = 63344;
	#10 counter$count = 63345;
	#10 counter$count = 63346;
	#10 counter$count = 63347;
	#10 counter$count = 63348;
	#10 counter$count = 63349;
	#10 counter$count = 63350;
	#10 counter$count = 63351;
	#10 counter$count = 63352;
	#10 counter$count = 63353;
	#10 counter$count = 63354;
	#10 counter$count = 63355;
	#10 counter$count = 63356;
	#10 counter$count = 63357;
	#10 counter$count = 63358;
	#10 counter$count = 63359;
	#10 counter$count = 63360;
	#10 counter$count = 63361;
	#10 counter$count = 63362;
	#10 counter$count = 63363;
	#10 counter$count = 63364;
	#10 counter$count = 63365;
	#10 counter$count = 63366;
	#10 counter$count = 63367;
	#10 counter$count = 63368;
	#10 counter$count = 63369;
	#10 counter$count = 63370;
	#10 counter$count = 63371;
	#10 counter$count = 63372;
	#10 counter$count = 63373;
	#10 counter$count = 63374;
	#10 counter$count = 63375;
	#10 counter$count = 63376;
	#10 counter$count = 63377;
	#10 counter$count = 63378;
	#10 counter$count = 63379;
	#10 counter$count = 63380;
	#10 counter$count = 63381;
	#10 counter$count = 63382;
	#10 counter$count = 63383;
	#10 counter$count = 63384;
	#10 counter$count = 63385;
	#10 counter$count = 63386;
	#10 counter$count = 63387;
	#10 counter$count = 63388;
	#10 counter$count = 63389;
	#10 counter$count = 63390;
	#10 counter$count = 63391;
	#10 counter$count = 63392;
	#10 counter$count = 63393;
	#10 counter$count = 63394;
	#10 counter$count = 63395;
	#10 counter$count = 63396;
	#10 counter$count = 63397;
	#10 counter$count = 63398;
	#10 counter$count = 63399;
	#10 counter$count = 63400;
	#10 counter$count = 63401;
	#10 counter$count = 63402;
	#10 counter$count = 63403;
	#10 counter$count = 63404;
	#10 counter$count = 63405;
	#10 counter$count = 63406;
	#10 counter$count = 63407;
	#10 counter$count = 63408;
	#10 counter$count = 63409;
	#10 counter$count = 63410;
	#10 counter$count = 63411;
	#10 counter$count = 63412;
	#10 counter$count = 63413;
	#10 counter$count = 63414;
	#10 counter$count = 63415;
	#10 counter$count = 63416;
	#10 counter$count = 63417;
	#10 counter$count = 63418;
	#10 counter$count = 63419;
	#10 counter$count = 63420;
	#10 counter$count = 63421;
	#10 counter$count = 63422;
	#10 counter$count = 63423;
	#10 counter$count = 63424;
	#10 counter$count = 63425;
	#10 counter$count = 63426;
	#10 counter$count = 63427;
	#10 counter$count = 63428;
	#10 counter$count = 63429;
	#10 counter$count = 63430;
	#10 counter$count = 63431;
	#10 counter$count = 63432;
	#10 counter$count = 63433;
	#10 counter$count = 63434;
	#10 counter$count = 63435;
	#10 counter$count = 63436;
	#10 counter$count = 63437;
	#10 counter$count = 63438;
	#10 counter$count = 63439;
	#10 counter$count = 63440;
	#10 counter$count = 63441;
	#10 counter$count = 63442;
	#10 counter$count = 63443;
	#10 counter$count = 63444;
	#10 counter$count = 63445;
	#10 counter$count = 63446;
	#10 counter$count = 63447;
	#10 counter$count = 63448;
	#10 counter$count = 63449;
	#10 counter$count = 63450;
	#10 counter$count = 63451;
	#10 counter$count = 63452;
	#10 counter$count = 63453;
	#10 counter$count = 63454;
	#10 counter$count = 63455;
	#10 counter$count = 63456;
	#10 counter$count = 63457;
	#10 counter$count = 63458;
	#10 counter$count = 63459;
	#10 counter$count = 63460;
	#10 counter$count = 63461;
	#10 counter$count = 63462;
	#10 counter$count = 63463;
	#10 counter$count = 63464;
	#10 counter$count = 63465;
	#10 counter$count = 63466;
	#10 counter$count = 63467;
	#10 counter$count = 63468;
	#10 counter$count = 63469;
	#10 counter$count = 63470;
	#10 counter$count = 63471;
	#10 counter$count = 63472;
	#10 counter$count = 63473;
	#10 counter$count = 63474;
	#10 counter$count = 63475;
	#10 counter$count = 63476;
	#10 counter$count = 63477;
	#10 counter$count = 63478;
	#10 counter$count = 63479;
	#10 counter$count = 63480;
	#10 counter$count = 63481;
	#10 counter$count = 63482;
	#10 counter$count = 63483;
	#10 counter$count = 63484;
	#10 counter$count = 63485;
	#10 counter$count = 63486;
	#10 counter$count = 63487;
	#10 counter$count = 63488;
	#10 counter$count = 63489;
	#10 counter$count = 63490;
	#10 counter$count = 63491;
	#10 counter$count = 63492;
	#10 counter$count = 63493;
	#10 counter$count = 63494;
	#10 counter$count = 63495;
	#10 counter$count = 63496;
	#10 counter$count = 63497;
	#10 counter$count = 63498;
	#10 counter$count = 63499;
	#10 counter$count = 63500;
	#10 counter$count = 63501;
	#10 counter$count = 63502;
	#10 counter$count = 63503;
	#10 counter$count = 63504;
	#10 counter$count = 63505;
	#10 counter$count = 63506;
	#10 counter$count = 63507;
	#10 counter$count = 63508;
	#10 counter$count = 63509;
	#10 counter$count = 63510;
	#10 counter$count = 63511;
	#10 counter$count = 63512;
	#10 counter$count = 63513;
	#10 counter$count = 63514;
	#10 counter$count = 63515;
	#10 counter$count = 63516;
	#10 counter$count = 63517;
	#10 counter$count = 63518;
	#10 counter$count = 63519;
	#10 counter$count = 63520;
	#10 counter$count = 63521;
	#10 counter$count = 63522;
	#10 counter$count = 63523;
	#10 counter$count = 63524;
	#10 counter$count = 63525;
	#10 counter$count = 63526;
	#10 counter$count = 63527;
	#10 counter$count = 63528;
	#10 counter$count = 63529;
	#10 counter$count = 63530;
	#10 counter$count = 63531;
	#10 counter$count = 63532;
	#10 counter$count = 63533;
	#10 counter$count = 63534;
	#10 counter$count = 63535;
	#10 counter$count = 63536;
	#10 counter$count = 63537;
	#10 counter$count = 63538;
	#10 counter$count = 63539;
	#10 counter$count = 63540;
	#10 counter$count = 63541;
	#10 counter$count = 63542;
	#10 counter$count = 63543;
	#10 counter$count = 63544;
	#10 counter$count = 63545;
	#10 counter$count = 63546;
	#10 counter$count = 63547;
	#10 counter$count = 63548;
	#10 counter$count = 63549;
	#10 counter$count = 63550;
	#10 counter$count = 63551;
	#10 counter$count = 63552;
	#10 counter$count = 63553;
	#10 counter$count = 63554;
	#10 counter$count = 63555;
	#10 counter$count = 63556;
	#10 counter$count = 63557;
	#10 counter$count = 63558;
	#10 counter$count = 63559;
	#10 counter$count = 63560;
	#10 counter$count = 63561;
	#10 counter$count = 63562;
	#10 counter$count = 63563;
	#10 counter$count = 63564;
	#10 counter$count = 63565;
	#10 counter$count = 63566;
	#10 counter$count = 63567;
	#10 counter$count = 63568;
	#10 counter$count = 63569;
	#10 counter$count = 63570;
	#10 counter$count = 63571;
	#10 counter$count = 63572;
	#10 counter$count = 63573;
	#10 counter$count = 63574;
	#10 counter$count = 63575;
	#10 counter$count = 63576;
	#10 counter$count = 63577;
	#10 counter$count = 63578;
	#10 counter$count = 63579;
	#10 counter$count = 63580;
	#10 counter$count = 63581;
	#10 counter$count = 63582;
	#10 counter$count = 63583;
	#10 counter$count = 63584;
	#10 counter$count = 63585;
	#10 counter$count = 63586;
	#10 counter$count = 63587;
	#10 counter$count = 63588;
	#10 counter$count = 63589;
	#10 counter$count = 63590;
	#10 counter$count = 63591;
	#10 counter$count = 63592;
	#10 counter$count = 63593;
	#10 counter$count = 63594;
	#10 counter$count = 63595;
	#10 counter$count = 63596;
	#10 counter$count = 63597;
	#10 counter$count = 63598;
	#10 counter$count = 63599;
	#10 counter$count = 63600;
	#10 counter$count = 63601;
	#10 counter$count = 63602;
	#10 counter$count = 63603;
	#10 counter$count = 63604;
	#10 counter$count = 63605;
	#10 counter$count = 63606;
	#10 counter$count = 63607;
	#10 counter$count = 63608;
	#10 counter$count = 63609;
	#10 counter$count = 63610;
	#10 counter$count = 63611;
	#10 counter$count = 63612;
	#10 counter$count = 63613;
	#10 counter$count = 63614;
	#10 counter$count = 63615;
	#10 counter$count = 63616;
	#10 counter$count = 63617;
	#10 counter$count = 63618;
	#10 counter$count = 63619;
	#10 counter$count = 63620;
	#10 counter$count = 63621;
	#10 counter$count = 63622;
	#10 counter$count = 63623;
	#10 counter$count = 63624;
	#10 counter$count = 63625;
	#10 counter$count = 63626;
	#10 counter$count = 63627;
	#10 counter$count = 63628;
	#10 counter$count = 63629;
	#10 counter$count = 63630;
	#10 counter$count = 63631;
	#10 counter$count = 63632;
	#10 counter$count = 63633;
	#10 counter$count = 63634;
	#10 counter$count = 63635;
	#10 counter$count = 63636;
	#10 counter$count = 63637;
	#10 counter$count = 63638;
	#10 counter$count = 63639;
	#10 counter$count = 63640;
	#10 counter$count = 63641;
	#10 counter$count = 63642;
	#10 counter$count = 63643;
	#10 counter$count = 63644;
	#10 counter$count = 63645;
	#10 counter$count = 63646;
	#10 counter$count = 63647;
	#10 counter$count = 63648;
	#10 counter$count = 63649;
	#10 counter$count = 63650;
	#10 counter$count = 63651;
	#10 counter$count = 63652;
	#10 counter$count = 63653;
	#10 counter$count = 63654;
	#10 counter$count = 63655;
	#10 counter$count = 63656;
	#10 counter$count = 63657;
	#10 counter$count = 63658;
	#10 counter$count = 63659;
	#10 counter$count = 63660;
	#10 counter$count = 63661;
	#10 counter$count = 63662;
	#10 counter$count = 63663;
	#10 counter$count = 63664;
	#10 counter$count = 63665;
	#10 counter$count = 63666;
	#10 counter$count = 63667;
	#10 counter$count = 63668;
	#10 counter$count = 63669;
	#10 counter$count = 63670;
	#10 counter$count = 63671;
	#10 counter$count = 63672;
	#10 counter$count = 63673;
	#10 counter$count = 63674;
	#10 counter$count = 63675;
	#10 counter$count = 63676;
	#10 counter$count = 63677;
	#10 counter$count = 63678;
	#10 counter$count = 63679;
	#10 counter$count = 63680;
	#10 counter$count = 63681;
	#10 counter$count = 63682;
	#10 counter$count = 63683;
	#10 counter$count = 63684;
	#10 counter$count = 63685;
	#10 counter$count = 63686;
	#10 counter$count = 63687;
	#10 counter$count = 63688;
	#10 counter$count = 63689;
	#10 counter$count = 63690;
	#10 counter$count = 63691;
	#10 counter$count = 63692;
	#10 counter$count = 63693;
	#10 counter$count = 63694;
	#10 counter$count = 63695;
	#10 counter$count = 63696;
	#10 counter$count = 63697;
	#10 counter$count = 63698;
	#10 counter$count = 63699;
	#10 counter$count = 63700;
	#10 counter$count = 63701;
	#10 counter$count = 63702;
	#10 counter$count = 63703;
	#10 counter$count = 63704;
	#10 counter$count = 63705;
	#10 counter$count = 63706;
	#10 counter$count = 63707;
	#10 counter$count = 63708;
	#10 counter$count = 63709;
	#10 counter$count = 63710;
	#10 counter$count = 63711;
	#10 counter$count = 63712;
	#10 counter$count = 63713;
	#10 counter$count = 63714;
	#10 counter$count = 63715;
	#10 counter$count = 63716;
	#10 counter$count = 63717;
	#10 counter$count = 63718;
	#10 counter$count = 63719;
	#10 counter$count = 63720;
	#10 counter$count = 63721;
	#10 counter$count = 63722;
	#10 counter$count = 63723;
	#10 counter$count = 63724;
	#10 counter$count = 63725;
	#10 counter$count = 63726;
	#10 counter$count = 63727;
	#10 counter$count = 63728;
	#10 counter$count = 63729;
	#10 counter$count = 63730;
	#10 counter$count = 63731;
	#10 counter$count = 63732;
	#10 counter$count = 63733;
	#10 counter$count = 63734;
	#10 counter$count = 63735;
	#10 counter$count = 63736;
	#10 counter$count = 63737;
	#10 counter$count = 63738;
	#10 counter$count = 63739;
	#10 counter$count = 63740;
	#10 counter$count = 63741;
	#10 counter$count = 63742;
	#10 counter$count = 63743;
	#10 counter$count = 63744;
	#10 counter$count = 63745;
	#10 counter$count = 63746;
	#10 counter$count = 63747;
	#10 counter$count = 63748;
	#10 counter$count = 63749;
	#10 counter$count = 63750;
	#10 counter$count = 63751;
	#10 counter$count = 63752;
	#10 counter$count = 63753;
	#10 counter$count = 63754;
	#10 counter$count = 63755;
	#10 counter$count = 63756;
	#10 counter$count = 63757;
	#10 counter$count = 63758;
	#10 counter$count = 63759;
	#10 counter$count = 63760;
	#10 counter$count = 63761;
	#10 counter$count = 63762;
	#10 counter$count = 63763;
	#10 counter$count = 63764;
	#10 counter$count = 63765;
	#10 counter$count = 63766;
	#10 counter$count = 63767;
	#10 counter$count = 63768;
	#10 counter$count = 63769;
	#10 counter$count = 63770;
	#10 counter$count = 63771;
	#10 counter$count = 63772;
	#10 counter$count = 63773;
	#10 counter$count = 63774;
	#10 counter$count = 63775;
	#10 counter$count = 63776;
	#10 counter$count = 63777;
	#10 counter$count = 63778;
	#10 counter$count = 63779;
	#10 counter$count = 63780;
	#10 counter$count = 63781;
	#10 counter$count = 63782;
	#10 counter$count = 63783;
	#10 counter$count = 63784;
	#10 counter$count = 63785;
	#10 counter$count = 63786;
	#10 counter$count = 63787;
	#10 counter$count = 63788;
	#10 counter$count = 63789;
	#10 counter$count = 63790;
	#10 counter$count = 63791;
	#10 counter$count = 63792;
	#10 counter$count = 63793;
	#10 counter$count = 63794;
	#10 counter$count = 63795;
	#10 counter$count = 63796;
	#10 counter$count = 63797;
	#10 counter$count = 63798;
	#10 counter$count = 63799;
	#10 counter$count = 63800;
	#10 counter$count = 63801;
	#10 counter$count = 63802;
	#10 counter$count = 63803;
	#10 counter$count = 63804;
	#10 counter$count = 63805;
	#10 counter$count = 63806;
	#10 counter$count = 63807;
	#10 counter$count = 63808;
	#10 counter$count = 63809;
	#10 counter$count = 63810;
	#10 counter$count = 63811;
	#10 counter$count = 63812;
	#10 counter$count = 63813;
	#10 counter$count = 63814;
	#10 counter$count = 63815;
	#10 counter$count = 63816;
	#10 counter$count = 63817;
	#10 counter$count = 63818;
	#10 counter$count = 63819;
	#10 counter$count = 63820;
	#10 counter$count = 63821;
	#10 counter$count = 63822;
	#10 counter$count = 63823;
	#10 counter$count = 63824;
	#10 counter$count = 63825;
	#10 counter$count = 63826;
	#10 counter$count = 63827;
	#10 counter$count = 63828;
	#10 counter$count = 63829;
	#10 counter$count = 63830;
	#10 counter$count = 63831;
	#10 counter$count = 63832;
	#10 counter$count = 63833;
	#10 counter$count = 63834;
	#10 counter$count = 63835;
	#10 counter$count = 63836;
	#10 counter$count = 63837;
	#10 counter$count = 63838;
	#10 counter$count = 63839;
	#10 counter$count = 63840;
	#10 counter$count = 63841;
	#10 counter$count = 63842;
	#10 counter$count = 63843;
	#10 counter$count = 63844;
	#10 counter$count = 63845;
	#10 counter$count = 63846;
	#10 counter$count = 63847;
	#10 counter$count = 63848;
	#10 counter$count = 63849;
	#10 counter$count = 63850;
	#10 counter$count = 63851;
	#10 counter$count = 63852;
	#10 counter$count = 63853;
	#10 counter$count = 63854;
	#10 counter$count = 63855;
	#10 counter$count = 63856;
	#10 counter$count = 63857;
	#10 counter$count = 63858;
	#10 counter$count = 63859;
	#10 counter$count = 63860;
	#10 counter$count = 63861;
	#10 counter$count = 63862;
	#10 counter$count = 63863;
	#10 counter$count = 63864;
	#10 counter$count = 63865;
	#10 counter$count = 63866;
	#10 counter$count = 63867;
	#10 counter$count = 63868;
	#10 counter$count = 63869;
	#10 counter$count = 63870;
	#10 counter$count = 63871;
	#10 counter$count = 63872;
	#10 counter$count = 63873;
	#10 counter$count = 63874;
	#10 counter$count = 63875;
	#10 counter$count = 63876;
	#10 counter$count = 63877;
	#10 counter$count = 63878;
	#10 counter$count = 63879;
	#10 counter$count = 63880;
	#10 counter$count = 63881;
	#10 counter$count = 63882;
	#10 counter$count = 63883;
	#10 counter$count = 63884;
	#10 counter$count = 63885;
	#10 counter$count = 63886;
	#10 counter$count = 63887;
	#10 counter$count = 63888;
	#10 counter$count = 63889;
	#10 counter$count = 63890;
	#10 counter$count = 63891;
	#10 counter$count = 63892;
	#10 counter$count = 63893;
	#10 counter$count = 63894;
	#10 counter$count = 63895;
	#10 counter$count = 63896;
	#10 counter$count = 63897;
	#10 counter$count = 63898;
	#10 counter$count = 63899;
	#10 counter$count = 63900;
	#10 counter$count = 63901;
	#10 counter$count = 63902;
	#10 counter$count = 63903;
	#10 counter$count = 63904;
	#10 counter$count = 63905;
	#10 counter$count = 63906;
	#10 counter$count = 63907;
	#10 counter$count = 63908;
	#10 counter$count = 63909;
	#10 counter$count = 63910;
	#10 counter$count = 63911;
	#10 counter$count = 63912;
	#10 counter$count = 63913;
	#10 counter$count = 63914;
	#10 counter$count = 63915;
	#10 counter$count = 63916;
	#10 counter$count = 63917;
	#10 counter$count = 63918;
	#10 counter$count = 63919;
	#10 counter$count = 63920;
	#10 counter$count = 63921;
	#10 counter$count = 63922;
	#10 counter$count = 63923;
	#10 counter$count = 63924;
	#10 counter$count = 63925;
	#10 counter$count = 63926;
	#10 counter$count = 63927;
	#10 counter$count = 63928;
	#10 counter$count = 63929;
	#10 counter$count = 63930;
	#10 counter$count = 63931;
	#10 counter$count = 63932;
	#10 counter$count = 63933;
	#10 counter$count = 63934;
	#10 counter$count = 63935;
	#10 counter$count = 63936;
	#10 counter$count = 63937;
	#10 counter$count = 63938;
	#10 counter$count = 63939;
	#10 counter$count = 63940;
	#10 counter$count = 63941;
	#10 counter$count = 63942;
	#10 counter$count = 63943;
	#10 counter$count = 63944;
	#10 counter$count = 63945;
	#10 counter$count = 63946;
	#10 counter$count = 63947;
	#10 counter$count = 63948;
	#10 counter$count = 63949;
	#10 counter$count = 63950;
	#10 counter$count = 63951;
	#10 counter$count = 63952;
	#10 counter$count = 63953;
	#10 counter$count = 63954;
	#10 counter$count = 63955;
	#10 counter$count = 63956;
	#10 counter$count = 63957;
	#10 counter$count = 63958;
	#10 counter$count = 63959;
	#10 counter$count = 63960;
	#10 counter$count = 63961;
	#10 counter$count = 63962;
	#10 counter$count = 63963;
	#10 counter$count = 63964;
	#10 counter$count = 63965;
	#10 counter$count = 63966;
	#10 counter$count = 63967;
	#10 counter$count = 63968;
	#10 counter$count = 63969;
	#10 counter$count = 63970;
	#10 counter$count = 63971;
	#10 counter$count = 63972;
	#10 counter$count = 63973;
	#10 counter$count = 63974;
	#10 counter$count = 63975;
	#10 counter$count = 63976;
	#10 counter$count = 63977;
	#10 counter$count = 63978;
	#10 counter$count = 63979;
	#10 counter$count = 63980;
	#10 counter$count = 63981;
	#10 counter$count = 63982;
	#10 counter$count = 63983;
	#10 counter$count = 63984;
	#10 counter$count = 63985;
	#10 counter$count = 63986;
	#10 counter$count = 63987;
	#10 counter$count = 63988;
	#10 counter$count = 63989;
	#10 counter$count = 63990;
	#10 counter$count = 63991;
	#10 counter$count = 63992;
	#10 counter$count = 63993;
	#10 counter$count = 63994;
	#10 counter$count = 63995;
	#10 counter$count = 63996;
	#10 counter$count = 63997;
	#10 counter$count = 63998;
	#10 counter$count = 63999;
	#10 counter$count = 64000;
	#10 counter$count = 64001;
	#10 counter$count = 64002;
	#10 counter$count = 64003;
	#10 counter$count = 64004;
	#10 counter$count = 64005;
	#10 counter$count = 64006;
	#10 counter$count = 64007;
	#10 counter$count = 64008;
	#10 counter$count = 64009;
	#10 counter$count = 64010;
	#10 counter$count = 64011;
	#10 counter$count = 64012;
	#10 counter$count = 64013;
	#10 counter$count = 64014;
	#10 counter$count = 64015;
	#10 counter$count = 64016;
	#10 counter$count = 64017;
	#10 counter$count = 64018;
	#10 counter$count = 64019;
	#10 counter$count = 64020;
	#10 counter$count = 64021;
	#10 counter$count = 64022;
	#10 counter$count = 64023;
	#10 counter$count = 64024;
	#10 counter$count = 64025;
	#10 counter$count = 64026;
	#10 counter$count = 64027;
	#10 counter$count = 64028;
	#10 counter$count = 64029;
	#10 counter$count = 64030;
	#10 counter$count = 64031;
	#10 counter$count = 64032;
	#10 counter$count = 64033;
	#10 counter$count = 64034;
	#10 counter$count = 64035;
	#10 counter$count = 64036;
	#10 counter$count = 64037;
	#10 counter$count = 64038;
	#10 counter$count = 64039;
	#10 counter$count = 64040;
	#10 counter$count = 64041;
	#10 counter$count = 64042;
	#10 counter$count = 64043;
	#10 counter$count = 64044;
	#10 counter$count = 64045;
	#10 counter$count = 64046;
	#10 counter$count = 64047;
	#10 counter$count = 64048;
	#10 counter$count = 64049;
	#10 counter$count = 64050;
	#10 counter$count = 64051;
	#10 counter$count = 64052;
	#10 counter$count = 64053;
	#10 counter$count = 64054;
	#10 counter$count = 64055;
	#10 counter$count = 64056;
	#10 counter$count = 64057;
	#10 counter$count = 64058;
	#10 counter$count = 64059;
	#10 counter$count = 64060;
	#10 counter$count = 64061;
	#10 counter$count = 64062;
	#10 counter$count = 64063;
	#10 counter$count = 64064;
	#10 counter$count = 64065;
	#10 counter$count = 64066;
	#10 counter$count = 64067;
	#10 counter$count = 64068;
	#10 counter$count = 64069;
	#10 counter$count = 64070;
	#10 counter$count = 64071;
	#10 counter$count = 64072;
	#10 counter$count = 64073;
	#10 counter$count = 64074;
	#10 counter$count = 64075;
	#10 counter$count = 64076;
	#10 counter$count = 64077;
	#10 counter$count = 64078;
	#10 counter$count = 64079;
	#10 counter$count = 64080;
	#10 counter$count = 64081;
	#10 counter$count = 64082;
	#10 counter$count = 64083;
	#10 counter$count = 64084;
	#10 counter$count = 64085;
	#10 counter$count = 64086;
	#10 counter$count = 64087;
	#10 counter$count = 64088;
	#10 counter$count = 64089;
	#10 counter$count = 64090;
	#10 counter$count = 64091;
	#10 counter$count = 64092;
	#10 counter$count = 64093;
	#10 counter$count = 64094;
	#10 counter$count = 64095;
	#10 counter$count = 64096;
	#10 counter$count = 64097;
	#10 counter$count = 64098;
	#10 counter$count = 64099;
	#10 counter$count = 64100;
	#10 counter$count = 64101;
	#10 counter$count = 64102;
	#10 counter$count = 64103;
	#10 counter$count = 64104;
	#10 counter$count = 64105;
	#10 counter$count = 64106;
	#10 counter$count = 64107;
	#10 counter$count = 64108;
	#10 counter$count = 64109;
	#10 counter$count = 64110;
	#10 counter$count = 64111;
	#10 counter$count = 64112;
	#10 counter$count = 64113;
	#10 counter$count = 64114;
	#10 counter$count = 64115;
	#10 counter$count = 64116;
	#10 counter$count = 64117;
	#10 counter$count = 64118;
	#10 counter$count = 64119;
	#10 counter$count = 64120;
	#10 counter$count = 64121;
	#10 counter$count = 64122;
	#10 counter$count = 64123;
	#10 counter$count = 64124;
	#10 counter$count = 64125;
	#10 counter$count = 64126;
	#10 counter$count = 64127;
	#10 counter$count = 64128;
	#10 counter$count = 64129;
	#10 counter$count = 64130;
	#10 counter$count = 64131;
	#10 counter$count = 64132;
	#10 counter$count = 64133;
	#10 counter$count = 64134;
	#10 counter$count = 64135;
	#10 counter$count = 64136;
	#10 counter$count = 64137;
	#10 counter$count = 64138;
	#10 counter$count = 64139;
	#10 counter$count = 64140;
	#10 counter$count = 64141;
	#10 counter$count = 64142;
	#10 counter$count = 64143;
	#10 counter$count = 64144;
	#10 counter$count = 64145;
	#10 counter$count = 64146;
	#10 counter$count = 64147;
	#10 counter$count = 64148;
	#10 counter$count = 64149;
	#10 counter$count = 64150;
	#10 counter$count = 64151;
	#10 counter$count = 64152;
	#10 counter$count = 64153;
	#10 counter$count = 64154;
	#10 counter$count = 64155;
	#10 counter$count = 64156;
	#10 counter$count = 64157;
	#10 counter$count = 64158;
	#10 counter$count = 64159;
	#10 counter$count = 64160;
	#10 counter$count = 64161;
	#10 counter$count = 64162;
	#10 counter$count = 64163;
	#10 counter$count = 64164;
	#10 counter$count = 64165;
	#10 counter$count = 64166;
	#10 counter$count = 64167;
	#10 counter$count = 64168;
	#10 counter$count = 64169;
	#10 counter$count = 64170;
	#10 counter$count = 64171;
	#10 counter$count = 64172;
	#10 counter$count = 64173;
	#10 counter$count = 64174;
	#10 counter$count = 64175;
	#10 counter$count = 64176;
	#10 counter$count = 64177;
	#10 counter$count = 64178;
	#10 counter$count = 64179;
	#10 counter$count = 64180;
	#10 counter$count = 64181;
	#10 counter$count = 64182;
	#10 counter$count = 64183;
	#10 counter$count = 64184;
	#10 counter$count = 64185;
	#10 counter$count = 64186;
	#10 counter$count = 64187;
	#10 counter$count = 64188;
	#10 counter$count = 64189;
	#10 counter$count = 64190;
	#10 counter$count = 64191;
	#10 counter$count = 64192;
	#10 counter$count = 64193;
	#10 counter$count = 64194;
	#10 counter$count = 64195;
	#10 counter$count = 64196;
	#10 counter$count = 64197;
	#10 counter$count = 64198;
	#10 counter$count = 64199;
	#10 counter$count = 64200;
	#10 counter$count = 64201;
	#10 counter$count = 64202;
	#10 counter$count = 64203;
	#10 counter$count = 64204;
	#10 counter$count = 64205;
	#10 counter$count = 64206;
	#10 counter$count = 64207;
	#10 counter$count = 64208;
	#10 counter$count = 64209;
	#10 counter$count = 64210;
	#10 counter$count = 64211;
	#10 counter$count = 64212;
	#10 counter$count = 64213;
	#10 counter$count = 64214;
	#10 counter$count = 64215;
	#10 counter$count = 64216;
	#10 counter$count = 64217;
	#10 counter$count = 64218;
	#10 counter$count = 64219;
	#10 counter$count = 64220;
	#10 counter$count = 64221;
	#10 counter$count = 64222;
	#10 counter$count = 64223;
	#10 counter$count = 64224;
	#10 counter$count = 64225;
	#10 counter$count = 64226;
	#10 counter$count = 64227;
	#10 counter$count = 64228;
	#10 counter$count = 64229;
	#10 counter$count = 64230;
	#10 counter$count = 64231;
	#10 counter$count = 64232;
	#10 counter$count = 64233;
	#10 counter$count = 64234;
	#10 counter$count = 64235;
	#10 counter$count = 64236;
	#10 counter$count = 64237;
	#10 counter$count = 64238;
	#10 counter$count = 64239;
	#10 counter$count = 64240;
	#10 counter$count = 64241;
	#10 counter$count = 64242;
	#10 counter$count = 64243;
	#10 counter$count = 64244;
	#10 counter$count = 64245;
	#10 counter$count = 64246;
	#10 counter$count = 64247;
	#10 counter$count = 64248;
	#10 counter$count = 64249;
	#10 counter$count = 64250;
	#10 counter$count = 64251;
	#10 counter$count = 64252;
	#10 counter$count = 64253;
	#10 counter$count = 64254;
	#10 counter$count = 64255;
	#10 counter$count = 64256;
	#10 counter$count = 64257;
	#10 counter$count = 64258;
	#10 counter$count = 64259;
	#10 counter$count = 64260;
	#10 counter$count = 64261;
	#10 counter$count = 64262;
	#10 counter$count = 64263;
	#10 counter$count = 64264;
	#10 counter$count = 64265;
	#10 counter$count = 64266;
	#10 counter$count = 64267;
	#10 counter$count = 64268;
	#10 counter$count = 64269;
	#10 counter$count = 64270;
	#10 counter$count = 64271;
	#10 counter$count = 64272;
	#10 counter$count = 64273;
	#10 counter$count = 64274;
	#10 counter$count = 64275;
	#10 counter$count = 64276;
	#10 counter$count = 64277;
	#10 counter$count = 64278;
	#10 counter$count = 64279;
	#10 counter$count = 64280;
	#10 counter$count = 64281;
	#10 counter$count = 64282;
	#10 counter$count = 64283;
	#10 counter$count = 64284;
	#10 counter$count = 64285;
	#10 counter$count = 64286;
	#10 counter$count = 64287;
	#10 counter$count = 64288;
	#10 counter$count = 64289;
	#10 counter$count = 64290;
	#10 counter$count = 64291;
	#10 counter$count = 64292;
	#10 counter$count = 64293;
	#10 counter$count = 64294;
	#10 counter$count = 64295;
	#10 counter$count = 64296;
	#10 counter$count = 64297;
	#10 counter$count = 64298;
	#10 counter$count = 64299;
	#10 counter$count = 64300;
	#10 counter$count = 64301;
	#10 counter$count = 64302;
	#10 counter$count = 64303;
	#10 counter$count = 64304;
	#10 counter$count = 64305;
	#10 counter$count = 64306;
	#10 counter$count = 64307;
	#10 counter$count = 64308;
	#10 counter$count = 64309;
	#10 counter$count = 64310;
	#10 counter$count = 64311;
	#10 counter$count = 64312;
	#10 counter$count = 64313;
	#10 counter$count = 64314;
	#10 counter$count = 64315;
	#10 counter$count = 64316;
	#10 counter$count = 64317;
	#10 counter$count = 64318;
	#10 counter$count = 64319;
	#10 counter$count = 64320;
	#10 counter$count = 64321;
	#10 counter$count = 64322;
	#10 counter$count = 64323;
	#10 counter$count = 64324;
	#10 counter$count = 64325;
	#10 counter$count = 64326;
	#10 counter$count = 64327;
	#10 counter$count = 64328;
	#10 counter$count = 64329;
	#10 counter$count = 64330;
	#10 counter$count = 64331;
	#10 counter$count = 64332;
	#10 counter$count = 64333;
	#10 counter$count = 64334;
	#10 counter$count = 64335;
	#10 counter$count = 64336;
	#10 counter$count = 64337;
	#10 counter$count = 64338;
	#10 counter$count = 64339;
	#10 counter$count = 64340;
	#10 counter$count = 64341;
	#10 counter$count = 64342;
	#10 counter$count = 64343;
	#10 counter$count = 64344;
	#10 counter$count = 64345;
	#10 counter$count = 64346;
	#10 counter$count = 64347;
	#10 counter$count = 64348;
	#10 counter$count = 64349;
	#10 counter$count = 64350;
	#10 counter$count = 64351;
	#10 counter$count = 64352;
	#10 counter$count = 64353;
	#10 counter$count = 64354;
	#10 counter$count = 64355;
	#10 counter$count = 64356;
	#10 counter$count = 64357;
	#10 counter$count = 64358;
	#10 counter$count = 64359;
	#10 counter$count = 64360;
	#10 counter$count = 64361;
	#10 counter$count = 64362;
	#10 counter$count = 64363;
	#10 counter$count = 64364;
	#10 counter$count = 64365;
	#10 counter$count = 64366;
	#10 counter$count = 64367;
	#10 counter$count = 64368;
	#10 counter$count = 64369;
	#10 counter$count = 64370;
	#10 counter$count = 64371;
	#10 counter$count = 64372;
	#10 counter$count = 64373;
	#10 counter$count = 64374;
	#10 counter$count = 64375;
	#10 counter$count = 64376;
	#10 counter$count = 64377;
	#10 counter$count = 64378;
	#10 counter$count = 64379;
	#10 counter$count = 64380;
	#10 counter$count = 64381;
	#10 counter$count = 64382;
	#10 counter$count = 64383;
	#10 counter$count = 64384;
	#10 counter$count = 64385;
	#10 counter$count = 64386;
	#10 counter$count = 64387;
	#10 counter$count = 64388;
	#10 counter$count = 64389;
	#10 counter$count = 64390;
	#10 counter$count = 64391;
	#10 counter$count = 64392;
	#10 counter$count = 64393;
	#10 counter$count = 64394;
	#10 counter$count = 64395;
	#10 counter$count = 64396;
	#10 counter$count = 64397;
	#10 counter$count = 64398;
	#10 counter$count = 64399;
	#10 counter$count = 64400;
	#10 counter$count = 64401;
	#10 counter$count = 64402;
	#10 counter$count = 64403;
	#10 counter$count = 64404;
	#10 counter$count = 64405;
	#10 counter$count = 64406;
	#10 counter$count = 64407;
	#10 counter$count = 64408;
	#10 counter$count = 64409;
	#10 counter$count = 64410;
	#10 counter$count = 64411;
	#10 counter$count = 64412;
	#10 counter$count = 64413;
	#10 counter$count = 64414;
	#10 counter$count = 64415;
	#10 counter$count = 64416;
	#10 counter$count = 64417;
	#10 counter$count = 64418;
	#10 counter$count = 64419;
	#10 counter$count = 64420;
	#10 counter$count = 64421;
	#10 counter$count = 64422;
	#10 counter$count = 64423;
	#10 counter$count = 64424;
	#10 counter$count = 64425;
	#10 counter$count = 64426;
	#10 counter$count = 64427;
	#10 counter$count = 64428;
	#10 counter$count = 64429;
	#10 counter$count = 64430;
	#10 counter$count = 64431;
	#10 counter$count = 64432;
	#10 counter$count = 64433;
	#10 counter$count = 64434;
	#10 counter$count = 64435;
	#10 counter$count = 64436;
	#10 counter$count = 64437;
	#10 counter$count = 64438;
	#10 counter$count = 64439;
	#10 counter$count = 64440;
	#10 counter$count = 64441;
	#10 counter$count = 64442;
	#10 counter$count = 64443;
	#10 counter$count = 64444;
	#10 counter$count = 64445;
	#10 counter$count = 64446;
	#10 counter$count = 64447;
	#10 counter$count = 64448;
	#10 counter$count = 64449;
	#10 counter$count = 64450;
	#10 counter$count = 64451;
	#10 counter$count = 64452;
	#10 counter$count = 64453;
	#10 counter$count = 64454;
	#10 counter$count = 64455;
	#10 counter$count = 64456;
	#10 counter$count = 64457;
	#10 counter$count = 64458;
	#10 counter$count = 64459;
	#10 counter$count = 64460;
	#10 counter$count = 64461;
	#10 counter$count = 64462;
	#10 counter$count = 64463;
	#10 counter$count = 64464;
	#10 counter$count = 64465;
	#10 counter$count = 64466;
	#10 counter$count = 64467;
	#10 counter$count = 64468;
	#10 counter$count = 64469;
	#10 counter$count = 64470;
	#10 counter$count = 64471;
	#10 counter$count = 64472;
	#10 counter$count = 64473;
	#10 counter$count = 64474;
	#10 counter$count = 64475;
	#10 counter$count = 64476;
	#10 counter$count = 64477;
	#10 counter$count = 64478;
	#10 counter$count = 64479;
	#10 counter$count = 64480;
	#10 counter$count = 64481;
	#10 counter$count = 64482;
	#10 counter$count = 64483;
	#10 counter$count = 64484;
	#10 counter$count = 64485;
	#10 counter$count = 64486;
	#10 counter$count = 64487;
	#10 counter$count = 64488;
	#10 counter$count = 64489;
	#10 counter$count = 64490;
	#10 counter$count = 64491;
	#10 counter$count = 64492;
	#10 counter$count = 64493;
	#10 counter$count = 64494;
	#10 counter$count = 64495;
	#10 counter$count = 64496;
	#10 counter$count = 64497;
	#10 counter$count = 64498;
	#10 counter$count = 64499;
	#10 counter$count = 64500;
	#10 counter$count = 64501;
	#10 counter$count = 64502;
	#10 counter$count = 64503;
	#10 counter$count = 64504;
	#10 counter$count = 64505;
	#10 counter$count = 64506;
	#10 counter$count = 64507;
	#10 counter$count = 64508;
	#10 counter$count = 64509;
	#10 counter$count = 64510;
	#10 counter$count = 64511;
	#10 counter$count = 64512;
	#10 counter$count = 64513;
	#10 counter$count = 64514;
	#10 counter$count = 64515;
	#10 counter$count = 64516;
	#10 counter$count = 64517;
	#10 counter$count = 64518;
	#10 counter$count = 64519;
	#10 counter$count = 64520;
	#10 counter$count = 64521;
	#10 counter$count = 64522;
	#10 counter$count = 64523;
	#10 counter$count = 64524;
	#10 counter$count = 64525;
	#10 counter$count = 64526;
	#10 counter$count = 64527;
	#10 counter$count = 64528;
	#10 counter$count = 64529;
	#10 counter$count = 64530;
	#10 counter$count = 64531;
	#10 counter$count = 64532;
	#10 counter$count = 64533;
	#10 counter$count = 64534;
	#10 counter$count = 64535;
	#10 counter$count = 64536;
	#10 counter$count = 64537;
	#10 counter$count = 64538;
	#10 counter$count = 64539;
	#10 counter$count = 64540;
	#10 counter$count = 64541;
	#10 counter$count = 64542;
	#10 counter$count = 64543;
	#10 counter$count = 64544;
	#10 counter$count = 64545;
	#10 counter$count = 64546;
	#10 counter$count = 64547;
	#10 counter$count = 64548;
	#10 counter$count = 64549;
	#10 counter$count = 64550;
	#10 counter$count = 64551;
	#10 counter$count = 64552;
	#10 counter$count = 64553;
	#10 counter$count = 64554;
	#10 counter$count = 64555;
	#10 counter$count = 64556;
	#10 counter$count = 64557;
	#10 counter$count = 64558;
	#10 counter$count = 64559;
	#10 counter$count = 64560;
	#10 counter$count = 64561;
	#10 counter$count = 64562;
	#10 counter$count = 64563;
	#10 counter$count = 64564;
	#10 counter$count = 64565;
	#10 counter$count = 64566;
	#10 counter$count = 64567;
	#10 counter$count = 64568;
	#10 counter$count = 64569;
	#10 counter$count = 64570;
	#10 counter$count = 64571;
	#10 counter$count = 64572;
	#10 counter$count = 64573;
	#10 counter$count = 64574;
	#10 counter$count = 64575;
	#10 counter$count = 64576;
	#10 counter$count = 64577;
	#10 counter$count = 64578;
	#10 counter$count = 64579;
	#10 counter$count = 64580;
	#10 counter$count = 64581;
	#10 counter$count = 64582;
	#10 counter$count = 64583;
	#10 counter$count = 64584;
	#10 counter$count = 64585;
	#10 counter$count = 64586;
	#10 counter$count = 64587;
	#10 counter$count = 64588;
	#10 counter$count = 64589;
	#10 counter$count = 64590;
	#10 counter$count = 64591;
	#10 counter$count = 64592;
	#10 counter$count = 64593;
	#10 counter$count = 64594;
	#10 counter$count = 64595;
	#10 counter$count = 64596;
	#10 counter$count = 64597;
	#10 counter$count = 64598;
	#10 counter$count = 64599;
	#10 counter$count = 64600;
	#10 counter$count = 64601;
	#10 counter$count = 64602;
	#10 counter$count = 64603;
	#10 counter$count = 64604;
	#10 counter$count = 64605;
	#10 counter$count = 64606;
	#10 counter$count = 64607;
	#10 counter$count = 64608;
	#10 counter$count = 64609;
	#10 counter$count = 64610;
	#10 counter$count = 64611;
	#10 counter$count = 64612;
	#10 counter$count = 64613;
	#10 counter$count = 64614;
	#10 counter$count = 64615;
	#10 counter$count = 64616;
	#10 counter$count = 64617;
	#10 counter$count = 64618;
	#10 counter$count = 64619;
	#10 counter$count = 64620;
	#10 counter$count = 64621;
	#10 counter$count = 64622;
	#10 counter$count = 64623;
	#10 counter$count = 64624;
	#10 counter$count = 64625;
	#10 counter$count = 64626;
	#10 counter$count = 64627;
	#10 counter$count = 64628;
	#10 counter$count = 64629;
	#10 counter$count = 64630;
	#10 counter$count = 64631;
	#10 counter$count = 64632;
	#10 counter$count = 64633;
	#10 counter$count = 64634;
	#10 counter$count = 64635;
	#10 counter$count = 64636;
	#10 counter$count = 64637;
	#10 counter$count = 64638;
	#10 counter$count = 64639;
	#10 counter$count = 64640;
	#10 counter$count = 64641;
	#10 counter$count = 64642;
	#10 counter$count = 64643;
	#10 counter$count = 64644;
	#10 counter$count = 64645;
	#10 counter$count = 64646;
	#10 counter$count = 64647;
	#10 counter$count = 64648;
	#10 counter$count = 64649;
	#10 counter$count = 64650;
	#10 counter$count = 64651;
	#10 counter$count = 64652;
	#10 counter$count = 64653;
	#10 counter$count = 64654;
	#10 counter$count = 64655;
	#10 counter$count = 64656;
	#10 counter$count = 64657;
	#10 counter$count = 64658;
	#10 counter$count = 64659;
	#10 counter$count = 64660;
	#10 counter$count = 64661;
	#10 counter$count = 64662;
	#10 counter$count = 64663;
	#10 counter$count = 64664;
	#10 counter$count = 64665;
	#10 counter$count = 64666;
	#10 counter$count = 64667;
	#10 counter$count = 64668;
	#10 counter$count = 64669;
	#10 counter$count = 64670;
	#10 counter$count = 64671;
	#10 counter$count = 64672;
	#10 counter$count = 64673;
	#10 counter$count = 64674;
	#10 counter$count = 64675;
	#10 counter$count = 64676;
	#10 counter$count = 64677;
	#10 counter$count = 64678;
	#10 counter$count = 64679;
	#10 counter$count = 64680;
	#10 counter$count = 64681;
	#10 counter$count = 64682;
	#10 counter$count = 64683;
	#10 counter$count = 64684;
	#10 counter$count = 64685;
	#10 counter$count = 64686;
	#10 counter$count = 64687;
	#10 counter$count = 64688;
	#10 counter$count = 64689;
	#10 counter$count = 64690;
	#10 counter$count = 64691;
	#10 counter$count = 64692;
	#10 counter$count = 64693;
	#10 counter$count = 64694;
	#10 counter$count = 64695;
	#10 counter$count = 64696;
	#10 counter$count = 64697;
	#10 counter$count = 64698;
	#10 counter$count = 64699;
	#10 counter$count = 64700;
	#10 counter$count = 64701;
	#10 counter$count = 64702;
	#10 counter$count = 64703;
	#10 counter$count = 64704;
	#10 counter$count = 64705;
	#10 counter$count = 64706;
	#10 counter$count = 64707;
	#10 counter$count = 64708;
	#10 counter$count = 64709;
	#10 counter$count = 64710;
	#10 counter$count = 64711;
	#10 counter$count = 64712;
	#10 counter$count = 64713;
	#10 counter$count = 64714;
	#10 counter$count = 64715;
	#10 counter$count = 64716;
	#10 counter$count = 64717;
	#10 counter$count = 64718;
	#10 counter$count = 64719;
	#10 counter$count = 64720;
	#10 counter$count = 64721;
	#10 counter$count = 64722;
	#10 counter$count = 64723;
	#10 counter$count = 64724;
	#10 counter$count = 64725;
	#10 counter$count = 64726;
	#10 counter$count = 64727;
	#10 counter$count = 64728;
	#10 counter$count = 64729;
	#10 counter$count = 64730;
	#10 counter$count = 64731;
	#10 counter$count = 64732;
	#10 counter$count = 64733;
	#10 counter$count = 64734;
	#10 counter$count = 64735;
	#10 counter$count = 64736;
	#10 counter$count = 64737;
	#10 counter$count = 64738;
	#10 counter$count = 64739;
	#10 counter$count = 64740;
	#10 counter$count = 64741;
	#10 counter$count = 64742;
	#10 counter$count = 64743;
	#10 counter$count = 64744;
	#10 counter$count = 64745;
	#10 counter$count = 64746;
	#10 counter$count = 64747;
	#10 counter$count = 64748;
	#10 counter$count = 64749;
	#10 counter$count = 64750;
	#10 counter$count = 64751;
	#10 counter$count = 64752;
	#10 counter$count = 64753;
	#10 counter$count = 64754;
	#10 counter$count = 64755;
	#10 counter$count = 64756;
	#10 counter$count = 64757;
	#10 counter$count = 64758;
	#10 counter$count = 64759;
	#10 counter$count = 64760;
	#10 counter$count = 64761;
	#10 counter$count = 64762;
	#10 counter$count = 64763;
	#10 counter$count = 64764;
	#10 counter$count = 64765;
	#10 counter$count = 64766;
	#10 counter$count = 64767;
	#10 counter$count = 64768;
	#10 counter$count = 64769;
	#10 counter$count = 64770;
	#10 counter$count = 64771;
	#10 counter$count = 64772;
	#10 counter$count = 64773;
	#10 counter$count = 64774;
	#10 counter$count = 64775;
	#10 counter$count = 64776;
	#10 counter$count = 64777;
	#10 counter$count = 64778;
	#10 counter$count = 64779;
	#10 counter$count = 64780;
	#10 counter$count = 64781;
	#10 counter$count = 64782;
	#10 counter$count = 64783;
	#10 counter$count = 64784;
	#10 counter$count = 64785;
	#10 counter$count = 64786;
	#10 counter$count = 64787;
	#10 counter$count = 64788;
	#10 counter$count = 64789;
	#10 counter$count = 64790;
	#10 counter$count = 64791;
	#10 counter$count = 64792;
	#10 counter$count = 64793;
	#10 counter$count = 64794;
	#10 counter$count = 64795;
	#10 counter$count = 64796;
	#10 counter$count = 64797;
	#10 counter$count = 64798;
	#10 counter$count = 64799;
	#10 counter$count = 64800;
	#10 counter$count = 64801;
	#10 counter$count = 64802;
	#10 counter$count = 64803;
	#10 counter$count = 64804;
	#10 counter$count = 64805;
	#10 counter$count = 64806;
	#10 counter$count = 64807;
	#10 counter$count = 64808;
	#10 counter$count = 64809;
	#10 counter$count = 64810;
	#10 counter$count = 64811;
	#10 counter$count = 64812;
	#10 counter$count = 64813;
	#10 counter$count = 64814;
	#10 counter$count = 64815;
	#10 counter$count = 64816;
	#10 counter$count = 64817;
	#10 counter$count = 64818;
	#10 counter$count = 64819;
	#10 counter$count = 64820;
	#10 counter$count = 64821;
	#10 counter$count = 64822;
	#10 counter$count = 64823;
	#10 counter$count = 64824;
	#10 counter$count = 64825;
	#10 counter$count = 64826;
	#10 counter$count = 64827;
	#10 counter$count = 64828;
	#10 counter$count = 64829;
	#10 counter$count = 64830;
	#10 counter$count = 64831;
	#10 counter$count = 64832;
	#10 counter$count = 64833;
	#10 counter$count = 64834;
	#10 counter$count = 64835;
	#10 counter$count = 64836;
	#10 counter$count = 64837;
	#10 counter$count = 64838;
	#10 counter$count = 64839;
	#10 counter$count = 64840;
	#10 counter$count = 64841;
	#10 counter$count = 64842;
	#10 counter$count = 64843;
	#10 counter$count = 64844;
	#10 counter$count = 64845;
	#10 counter$count = 64846;
	#10 counter$count = 64847;
	#10 counter$count = 64848;
	#10 counter$count = 64849;
	#10 counter$count = 64850;
	#10 counter$count = 64851;
	#10 counter$count = 64852;
	#10 counter$count = 64853;
	#10 counter$count = 64854;
	#10 counter$count = 64855;
	#10 counter$count = 64856;
	#10 counter$count = 64857;
	#10 counter$count = 64858;
	#10 counter$count = 64859;
	#10 counter$count = 64860;
	#10 counter$count = 64861;
	#10 counter$count = 64862;
	#10 counter$count = 64863;
	#10 counter$count = 64864;
	#10 counter$count = 64865;
	#10 counter$count = 64866;
	#10 counter$count = 64867;
	#10 counter$count = 64868;
	#10 counter$count = 64869;
	#10 counter$count = 64870;
	#10 counter$count = 64871;
	#10 counter$count = 64872;
	#10 counter$count = 64873;
	#10 counter$count = 64874;
	#10 counter$count = 64875;
	#10 counter$count = 64876;
	#10 counter$count = 64877;
	#10 counter$count = 64878;
	#10 counter$count = 64879;
	#10 counter$count = 64880;
	#10 counter$count = 64881;
	#10 counter$count = 64882;
	#10 counter$count = 64883;
	#10 counter$count = 64884;
	#10 counter$count = 64885;
	#10 counter$count = 64886;
	#10 counter$count = 64887;
	#10 counter$count = 64888;
	#10 counter$count = 64889;
	#10 counter$count = 64890;
	#10 counter$count = 64891;
	#10 counter$count = 64892;
	#10 counter$count = 64893;
	#10 counter$count = 64894;
	#10 counter$count = 64895;
	#10 counter$count = 64896;
	#10 counter$count = 64897;
	#10 counter$count = 64898;
	#10 counter$count = 64899;
	#10 counter$count = 64900;
	#10 counter$count = 64901;
	#10 counter$count = 64902;
	#10 counter$count = 64903;
	#10 counter$count = 64904;
	#10 counter$count = 64905;
	#10 counter$count = 64906;
	#10 counter$count = 64907;
	#10 counter$count = 64908;
	#10 counter$count = 64909;
	#10 counter$count = 64910;
	#10 counter$count = 64911;
	#10 counter$count = 64912;
	#10 counter$count = 64913;
	#10 counter$count = 64914;
	#10 counter$count = 64915;
	#10 counter$count = 64916;
	#10 counter$count = 64917;
	#10 counter$count = 64918;
	#10 counter$count = 64919;
	#10 counter$count = 64920;
	#10 counter$count = 64921;
	#10 counter$count = 64922;
	#10 counter$count = 64923;
	#10 counter$count = 64924;
	#10 counter$count = 64925;
	#10 counter$count = 64926;
	#10 counter$count = 64927;
	#10 counter$count = 64928;
	#10 counter$count = 64929;
	#10 counter$count = 64930;
	#10 counter$count = 64931;
	#10 counter$count = 64932;
	#10 counter$count = 64933;
	#10 counter$count = 64934;
	#10 counter$count = 64935;
	#10 counter$count = 64936;
	#10 counter$count = 64937;
	#10 counter$count = 64938;
	#10 counter$count = 64939;
	#10 counter$count = 64940;
	#10 counter$count = 64941;
	#10 counter$count = 64942;
	#10 counter$count = 64943;
	#10 counter$count = 64944;
	#10 counter$count = 64945;
	#10 counter$count = 64946;
	#10 counter$count = 64947;
	#10 counter$count = 64948;
	#10 counter$count = 64949;
	#10 counter$count = 64950;
	#10 counter$count = 64951;
	#10 counter$count = 64952;
	#10 counter$count = 64953;
	#10 counter$count = 64954;
	#10 counter$count = 64955;
	#10 counter$count = 64956;
	#10 counter$count = 64957;
	#10 counter$count = 64958;
	#10 counter$count = 64959;
	#10 counter$count = 64960;
	#10 counter$count = 64961;
	#10 counter$count = 64962;
	#10 counter$count = 64963;
	#10 counter$count = 64964;
	#10 counter$count = 64965;
	#10 counter$count = 64966;
	#10 counter$count = 64967;
	#10 counter$count = 64968;
	#10 counter$count = 64969;
	#10 counter$count = 64970;
	#10 counter$count = 64971;
	#10 counter$count = 64972;
	#10 counter$count = 64973;
	#10 counter$count = 64974;
	#10 counter$count = 64975;
	#10 counter$count = 64976;
	#10 counter$count = 64977;
	#10 counter$count = 64978;
	#10 counter$count = 64979;
	#10 counter$count = 64980;
	#10 counter$count = 64981;
	#10 counter$count = 64982;
	#10 counter$count = 64983;
	#10 counter$count = 64984;
	#10 counter$count = 64985;
	#10 counter$count = 64986;
	#10 counter$count = 64987;
	#10 counter$count = 64988;
	#10 counter$count = 64989;
	#10 counter$count = 64990;
	#10 counter$count = 64991;
	#10 counter$count = 64992;
	#10 counter$count = 64993;
	#10 counter$count = 64994;
	#10 counter$count = 64995;
	#10 counter$count = 64996;
	#10 counter$count = 64997;
	#10 counter$count = 64998;
	#10 counter$count = 64999;
	#10 counter$count = 65000;
	#10 counter$count = 65001;
	#10 counter$count = 65002;
	#10 counter$count = 65003;
	#10 counter$count = 65004;
	#10 counter$count = 65005;
	#10 counter$count = 65006;
	#10 counter$count = 65007;
	#10 counter$count = 65008;
	#10 counter$count = 65009;
	#10 counter$count = 65010;
	#10 counter$count = 65011;
	#10 counter$count = 65012;
	#10 counter$count = 65013;
	#10 counter$count = 65014;
	#10 counter$count = 65015;
	#10 counter$count = 65016;
	#10 counter$count = 65017;
	#10 counter$count = 65018;
	#10 counter$count = 65019;
	#10 counter$count = 65020;
	#10 counter$count = 65021;
	#10 counter$count = 65022;
	#10 counter$count = 65023;
	#10 counter$count = 65024;
	#10 counter$count = 65025;
	#10 counter$count = 65026;
	#10 counter$count = 65027;
	#10 counter$count = 65028;
	#10 counter$count = 65029;
	#10 counter$count = 65030;
	#10 counter$count = 65031;
	#10 counter$count = 65032;
	#10 counter$count = 65033;
	#10 counter$count = 65034;
	#10 counter$count = 65035;
	#10 counter$count = 65036;
	#10 counter$count = 65037;
	#10 counter$count = 65038;
	#10 counter$count = 65039;
	#10 counter$count = 65040;
	#10 counter$count = 65041;
	#10 counter$count = 65042;
	#10 counter$count = 65043;
	#10 counter$count = 65044;
	#10 counter$count = 65045;
	#10 counter$count = 65046;
	#10 counter$count = 65047;
	#10 counter$count = 65048;
	#10 counter$count = 65049;
	#10 counter$count = 65050;
	#10 counter$count = 65051;
	#10 counter$count = 65052;
	#10 counter$count = 65053;
	#10 counter$count = 65054;
	#10 counter$count = 65055;
	#10 counter$count = 65056;
	#10 counter$count = 65057;
	#10 counter$count = 65058;
	#10 counter$count = 65059;
	#10 counter$count = 65060;
	#10 counter$count = 65061;
	#10 counter$count = 65062;
	#10 counter$count = 65063;
	#10 counter$count = 65064;
	#10 counter$count = 65065;
	#10 counter$count = 65066;
	#10 counter$count = 65067;
	#10 counter$count = 65068;
	#10 counter$count = 65069;
	#10 counter$count = 65070;
	#10 counter$count = 65071;
	#10 counter$count = 65072;
	#10 counter$count = 65073;
	#10 counter$count = 65074;
	#10 counter$count = 65075;
	#10 counter$count = 65076;
	#10 counter$count = 65077;
	#10 counter$count = 65078;
	#10 counter$count = 65079;
	#10 counter$count = 65080;
	#10 counter$count = 65081;
	#10 counter$count = 65082;
	#10 counter$count = 65083;
	#10 counter$count = 65084;
	#10 counter$count = 65085;
	#10 counter$count = 65086;
	#10 counter$count = 65087;
	#10 counter$count = 65088;
	#10 counter$count = 65089;
	#10 counter$count = 65090;
	#10 counter$count = 65091;
	#10 counter$count = 65092;
	#10 counter$count = 65093;
	#10 counter$count = 65094;
	#10 counter$count = 65095;
	#10 counter$count = 65096;
	#10 counter$count = 65097;
	#10 counter$count = 65098;
	#10 counter$count = 65099;
	#10 counter$count = 65100;
	#10 counter$count = 65101;
	#10 counter$count = 65102;
	#10 counter$count = 65103;
	#10 counter$count = 65104;
	#10 counter$count = 65105;
	#10 counter$count = 65106;
	#10 counter$count = 65107;
	#10 counter$count = 65108;
	#10 counter$count = 65109;
	#10 counter$count = 65110;
	#10 counter$count = 65111;
	#10 counter$count = 65112;
	#10 counter$count = 65113;
	#10 counter$count = 65114;
	#10 counter$count = 65115;
	#10 counter$count = 65116;
	#10 counter$count = 65117;
	#10 counter$count = 65118;
	#10 counter$count = 65119;
	#10 counter$count = 65120;
	#10 counter$count = 65121;
	#10 counter$count = 65122;
	#10 counter$count = 65123;
	#10 counter$count = 65124;
	#10 counter$count = 65125;
	#10 counter$count = 65126;
	#10 counter$count = 65127;
	#10 counter$count = 65128;
	#10 counter$count = 65129;
	#10 counter$count = 65130;
	#10 counter$count = 65131;
	#10 counter$count = 65132;
	#10 counter$count = 65133;
	#10 counter$count = 65134;
	#10 counter$count = 65135;
	#10 counter$count = 65136;
	#10 counter$count = 65137;
	#10 counter$count = 65138;
	#10 counter$count = 65139;
	#10 counter$count = 65140;
	#10 counter$count = 65141;
	#10 counter$count = 65142;
	#10 counter$count = 65143;
	#10 counter$count = 65144;
	#10 counter$count = 65145;
	#10 counter$count = 65146;
	#10 counter$count = 65147;
	#10 counter$count = 65148;
	#10 counter$count = 65149;
	#10 counter$count = 65150;
	#10 counter$count = 65151;
	#10 counter$count = 65152;
	#10 counter$count = 65153;
	#10 counter$count = 65154;
	#10 counter$count = 65155;
	#10 counter$count = 65156;
	#10 counter$count = 65157;
	#10 counter$count = 65158;
	#10 counter$count = 65159;
	#10 counter$count = 65160;
	#10 counter$count = 65161;
	#10 counter$count = 65162;
	#10 counter$count = 65163;
	#10 counter$count = 65164;
	#10 counter$count = 65165;
	#10 counter$count = 65166;
	#10 counter$count = 65167;
	#10 counter$count = 65168;
	#10 counter$count = 65169;
	#10 counter$count = 65170;
	#10 counter$count = 65171;
	#10 counter$count = 65172;
	#10 counter$count = 65173;
	#10 counter$count = 65174;
	#10 counter$count = 65175;
	#10 counter$count = 65176;
	#10 counter$count = 65177;
	#10 counter$count = 65178;
	#10 counter$count = 65179;
	#10 counter$count = 65180;
	#10 counter$count = 65181;
	#10 counter$count = 65182;
	#10 counter$count = 65183;
	#10 counter$count = 65184;
	#10 counter$count = 65185;
	#10 counter$count = 65186;
	#10 counter$count = 65187;
	#10 counter$count = 65188;
	#10 counter$count = 65189;
	#10 counter$count = 65190;
	#10 counter$count = 65191;
	#10 counter$count = 65192;
	#10 counter$count = 65193;
	#10 counter$count = 65194;
	#10 counter$count = 65195;
	#10 counter$count = 65196;
	#10 counter$count = 65197;
	#10 counter$count = 65198;
	#10 counter$count = 65199;
	#10 counter$count = 65200;
	#10 counter$count = 65201;
	#10 counter$count = 65202;
	#10 counter$count = 65203;
	#10 counter$count = 65204;
	#10 counter$count = 65205;
	#10 counter$count = 65206;
	#10 counter$count = 65207;
	#10 counter$count = 65208;
	#10 counter$count = 65209;
	#10 counter$count = 65210;
	#10 counter$count = 65211;
	#10 counter$count = 65212;
	#10 counter$count = 65213;
	#10 counter$count = 65214;
	#10 counter$count = 65215;
	#10 counter$count = 65216;
	#10 counter$count = 65217;
	#10 counter$count = 65218;
	#10 counter$count = 65219;
	#10 counter$count = 65220;
	#10 counter$count = 65221;
	#10 counter$count = 65222;
	#10 counter$count = 65223;
	#10 counter$count = 65224;
	#10 counter$count = 65225;
	#10 counter$count = 65226;
	#10 counter$count = 65227;
	#10 counter$count = 65228;
	#10 counter$count = 65229;
	#10 counter$count = 65230;
	#10 counter$count = 65231;
	#10 counter$count = 65232;
	#10 counter$count = 65233;
	#10 counter$count = 65234;
	#10 counter$count = 65235;
	#10 counter$count = 65236;
	#10 counter$count = 65237;
	#10 counter$count = 65238;
	#10 counter$count = 65239;
	#10 counter$count = 65240;
	#10 counter$count = 65241;
	#10 counter$count = 65242;
	#10 counter$count = 65243;
	#10 counter$count = 65244;
	#10 counter$count = 65245;
	#10 counter$count = 65246;
	#10 counter$count = 65247;
	#10 counter$count = 65248;
	#10 counter$count = 65249;
	#10 counter$count = 65250;
	#10 counter$count = 65251;
	#10 counter$count = 65252;
	#10 counter$count = 65253;
	#10 counter$count = 65254;
	#10 counter$count = 65255;
	#10 counter$count = 65256;
	#10 counter$count = 65257;
	#10 counter$count = 65258;
	#10 counter$count = 65259;
	#10 counter$count = 65260;
	#10 counter$count = 65261;
	#10 counter$count = 65262;
	#10 counter$count = 65263;
	#10 counter$count = 65264;
	#10 counter$count = 65265;
	#10 counter$count = 65266;
	#10 counter$count = 65267;
	#10 counter$count = 65268;
	#10 counter$count = 65269;
	#10 counter$count = 65270;
	#10 counter$count = 65271;
	#10 counter$count = 65272;
	#10 counter$count = 65273;
	#10 counter$count = 65274;
	#10 counter$count = 65275;
	#10 counter$count = 65276;
	#10 counter$count = 65277;
	#10 counter$count = 65278;
	#10 counter$count = 65279;
	#10 counter$count = 65280;
	#10 counter$count = 65281;
	#10 counter$count = 65282;
	#10 counter$count = 65283;
	#10 counter$count = 65284;
	#10 counter$count = 65285;
	#10 counter$count = 65286;
	#10 counter$count = 65287;
	#10 counter$count = 65288;
	#10 counter$count = 65289;
	#10 counter$count = 65290;
	#10 counter$count = 65291;
	#10 counter$count = 65292;
	#10 counter$count = 65293;
	#10 counter$count = 65294;
	#10 counter$count = 65295;
	#10 counter$count = 65296;
	#10 counter$count = 65297;
	#10 counter$count = 65298;
	#10 counter$count = 65299;
	#10 counter$count = 65300;
	#10 counter$count = 65301;
	#10 counter$count = 65302;
	#10 counter$count = 65303;
	#10 counter$count = 65304;
	#10 counter$count = 65305;
	#10 counter$count = 65306;
	#10 counter$count = 65307;
	#10 counter$count = 65308;
	#10 counter$count = 65309;
	#10 counter$count = 65310;
	#10 counter$count = 65311;
	#10 counter$count = 65312;
	#10 counter$count = 65313;
	#10 counter$count = 65314;
	#10 counter$count = 65315;
	#10 counter$count = 65316;
	#10 counter$count = 65317;
	#10 counter$count = 65318;
	#10 counter$count = 65319;
	#10 counter$count = 65320;
	#10 counter$count = 65321;
	#10 counter$count = 65322;
	#10 counter$count = 65323;
	#10 counter$count = 65324;
	#10 counter$count = 65325;
	#10 counter$count = 65326;
	#10 counter$count = 65327;
	#10 counter$count = 65328;
	#10 counter$count = 65329;
	#10 counter$count = 65330;
	#10 counter$count = 65331;
	#10 counter$count = 65332;
	#10 counter$count = 65333;
	#10 counter$count = 65334;
	#10 counter$count = 65335;
	#10 counter$count = 65336;
	#10 counter$count = 65337;
	#10 counter$count = 65338;
	#10 counter$count = 65339;
	#10 counter$count = 65340;
	#10 counter$count = 65341;
	#10 counter$count = 65342;
	#10 counter$count = 65343;
	#10 counter$count = 65344;
	#10 counter$count = 65345;
	#10 counter$count = 65346;
	#10 counter$count = 65347;
	#10 counter$count = 65348;
	#10 counter$count = 65349;
	#10 counter$count = 65350;
	#10 counter$count = 65351;
	#10 counter$count = 65352;
	#10 counter$count = 65353;
	#10 counter$count = 65354;
	#10 counter$count = 65355;
	#10 counter$count = 65356;
	#10 counter$count = 65357;
	#10 counter$count = 65358;
	#10 counter$count = 65359;
	#10 counter$count = 65360;
	#10 counter$count = 65361;
	#10 counter$count = 65362;
	#10 counter$count = 65363;
	#10 counter$count = 65364;
	#10 counter$count = 65365;
	#10 counter$count = 65366;
	#10 counter$count = 65367;
	#10 counter$count = 65368;
	#10 counter$count = 65369;
	#10 counter$count = 65370;
	#10 counter$count = 65371;
	#10 counter$count = 65372;
	#10 counter$count = 65373;
	#10 counter$count = 65374;
	#10 counter$count = 65375;
	#10 counter$count = 65376;
	#10 counter$count = 65377;
	#10 counter$count = 65378;
	#10 counter$count = 65379;
	#10 counter$count = 65380;
	#10 counter$count = 65381;
	#10 counter$count = 65382;
	#10 counter$count = 65383;
	#10 counter$count = 65384;
	#10 counter$count = 65385;
	#10 counter$count = 65386;
	#10 counter$count = 65387;
	#10 counter$count = 65388;
	#10 counter$count = 65389;
	#10 counter$count = 65390;
	#10 counter$count = 65391;
	#10 counter$count = 65392;
	#10 counter$count = 65393;
	#10 counter$count = 65394;
	#10 counter$count = 65395;
	#10 counter$count = 65396;
	#10 counter$count = 65397;
	#10 counter$count = 65398;
	#10 counter$count = 65399;
	#10 counter$count = 65400;
	#10 counter$count = 65401;
	#10 counter$count = 65402;
	#10 counter$count = 65403;
	#10 counter$count = 65404;
	#10 counter$count = 65405;
	#10 counter$count = 65406;
	#10 counter$count = 65407;
	#10 counter$count = 65408;
	#10 counter$count = 65409;
	#10 counter$count = 65410;
	#10 counter$count = 65411;
	#10 counter$count = 65412;
	#10 counter$count = 65413;
	#10 counter$count = 65414;
	#10 counter$count = 65415;
	#10 counter$count = 65416;
	#10 counter$count = 65417;
	#10 counter$count = 65418;
	#10 counter$count = 65419;
	#10 counter$count = 65420;
	#10 counter$count = 65421;
	#10 counter$count = 65422;
	#10 counter$count = 65423;
	#10 counter$count = 65424;
	#10 counter$count = 65425;
	#10 counter$count = 65426;
	#10 counter$count = 65427;
	#10 counter$count = 65428;
	#10 counter$count = 65429;
	#10 counter$count = 65430;
	#10 counter$count = 65431;
	#10 counter$count = 65432;
	#10 counter$count = 65433;
	#10 counter$count = 65434;
	#10 counter$count = 65435;
	#10 counter$count = 65436;
	#10 counter$count = 65437;
	#10 counter$count = 65438;
	#10 counter$count = 65439;
	#10 counter$count = 65440;
	#10 counter$count = 65441;
	#10 counter$count = 65442;
	#10 counter$count = 65443;
	#10 counter$count = 65444;
	#10 counter$count = 65445;
	#10 counter$count = 65446;
	#10 counter$count = 65447;
	#10 counter$count = 65448;
	#10 counter$count = 65449;
	#10 counter$count = 65450;
	#10 counter$count = 65451;
	#10 counter$count = 65452;
	#10 counter$count = 65453;
	#10 counter$count = 65454;
	#10 counter$count = 65455;
	#10 counter$count = 65456;
	#10 counter$count = 65457;
	#10 counter$count = 65458;
	#10 counter$count = 65459;
	#10 counter$count = 65460;
	#10 counter$count = 65461;
	#10 counter$count = 65462;
	#10 counter$count = 65463;
	#10 counter$count = 65464;
	#10 counter$count = 65465;
	#10 counter$count = 65466;
	#10 counter$count = 65467;
	#10 counter$count = 65468;
	#10 counter$count = 65469;
	#10 counter$count = 65470;
	#10 counter$count = 65471;
	#10 counter$count = 65472;
	#10 counter$count = 65473;
	#10 counter$count = 65474;
	#10 counter$count = 65475;
	#10 counter$count = 65476;
	#10 counter$count = 65477;
	#10 counter$count = 65478;
	#10 counter$count = 65479;
	#10 counter$count = 65480;
	#10 counter$count = 65481;
	#10 counter$count = 65482;
	#10 counter$count = 65483;
	#10 counter$count = 65484;
	#10 counter$count = 65485;
	#10 counter$count = 65486;
	#10 counter$count = 65487;
	#10 counter$count = 65488;
	#10 counter$count = 65489;
	#10 counter$count = 65490;
	#10 counter$count = 65491;
	#10 counter$count = 65492;
	#10 counter$count = 65493;
	#10 counter$count = 65494;
	#10 counter$count = 65495;
	#10 counter$count = 65496;
	#10 counter$count = 65497;
	#10 counter$count = 65498;
	#10 counter$count = 65499;
	#10 counter$count = 65500;
	#10 counter$count = 65501;
	#10 counter$count = 65502;
	#10 counter$count = 65503;
	#10 counter$count = 65504;
	#10 counter$count = 65505;
	#10 counter$count = 65506;
	#10 counter$count = 65507;
	#10 counter$count = 65508;
	#10 counter$count = 65509;
	#10 counter$count = 65510;
	#10 counter$count = 65511;
	#10 counter$count = 65512;
	#10 counter$count = 65513;
	#10 counter$count = 65514;
	#10 counter$count = 65515;
	#10 counter$count = 65516;
	#10 counter$count = 65517;
	#10 counter$count = 65518;
	#10 counter$count = 65519;
	#10 counter$count = 65520;
	#10 counter$count = 65521;
	#10 counter$count = 65522;
	#10 counter$count = 65523;
	#10 counter$count = 65524;
	#10 counter$count = 65525;
	#10 counter$count = 65526;
	#10 counter$count = 65527;
	#10 counter$count = 65528;
	#10 counter$count = 65529;
	#10 counter$count = 65530;
	#10 counter$count = 65531;
	#10 counter$count = 65532;
	#10 counter$count = 65533;
	#10 counter$count = 65534;
	#10 counter$count = 65535;
	#10 counter$count = 65536;
	#10 counter$count = 65537;
	#10 counter$count = 65538;
	#10 counter$count = 65539;
	#10 counter$count = 65540;
	#10 counter$count = 65541;
	#10 counter$count = 65542;
	#10 counter$count = 65543;
	#10 counter$count = 65544;
	#10 counter$count = 65545;
	#10 counter$count = 65546;
	#10 counter$count = 65547;
	#10 counter$count = 65548;
	#10 counter$count = 65549;
	#10 counter$count = 65550;
	#10 counter$count = 65551;
	#10 counter$count = 65552;
	#10 counter$count = 65553;
	#10 counter$count = 65554;
	#10 counter$count = 65555;
	#10 counter$count = 65556;
	#10 counter$count = 65557;
	#10 counter$count = 65558;
	#10 counter$count = 65559;
	#10 counter$count = 65560;
	#10 counter$count = 65561;
	#10 counter$count = 65562;
	#10 counter$count = 65563;
	#10 counter$count = 65564;
	#10 counter$count = 65565;
	#10 counter$count = 65566;
	#10 counter$count = 65567;
	#10 counter$count = 65568;
	#10 counter$count = 65569;
	#10 counter$count = 65570;
	#10 counter$count = 65571;
	#10 counter$count = 65572;
	#10 counter$count = 65573;
	#10 counter$count = 65574;
	#10 counter$count = 65575;
	#10 counter$count = 65576;
	#10 counter$count = 65577;
	#10 counter$count = 65578;
	#10 counter$count = 65579;
	#10 counter$count = 65580;
	#10 counter$count = 65581;
	#10 counter$count = 65582;
	#10 counter$count = 65583;
	#10 counter$count = 65584;
	#10 counter$count = 65585;
	#10 counter$count = 65586;
	#10 counter$count = 65587;
	#10 counter$count = 65588;
	#10 counter$count = 65589;
	#10 counter$count = 65590;
	#10 counter$count = 65591;
	#10 counter$count = 65592;
	#10 counter$count = 65593;
	#10 counter$count = 65594;
	#10 counter$count = 65595;
	#10 counter$count = 65596;
	#10 counter$count = 65597;
	#10 counter$count = 65598;
	#10 counter$count = 65599;
	#10 counter$count = 65600;
	#10 counter$count = 65601;
	#10 counter$count = 65602;
	#10 counter$count = 65603;
	#10 counter$count = 65604;
	#10 counter$count = 65605;
	#10 counter$count = 65606;
	#10 counter$count = 65607;
	#10 counter$count = 65608;
	#10 counter$count = 65609;
	#10 counter$count = 65610;
	#10 counter$count = 65611;
	#10 counter$count = 65612;
	#10 counter$count = 65613;
	#10 counter$count = 65614;
	#10 counter$count = 65615;
	#10 counter$count = 65616;
	#10 counter$count = 65617;
	#10 counter$count = 65618;
	#10 counter$count = 65619;
	#10 counter$count = 65620;
	#10 counter$count = 65621;
	#10 counter$count = 65622;
	#10 counter$count = 65623;
	#10 counter$count = 65624;
	#10 counter$count = 65625;
	#10 counter$count = 65626;
	#10 counter$count = 65627;
	#10 counter$count = 65628;
	#10 counter$count = 65629;
	#10 counter$count = 65630;
	#10 counter$count = 65631;
	#10 counter$count = 65632;
	#10 counter$count = 65633;
	#10 counter$count = 65634;
	#10 counter$count = 65635;
	#10 counter$count = 65636;
	#10 counter$count = 65637;
	#10 counter$count = 65638;
	#10 counter$count = 65639;
	#10 counter$count = 65640;
	#10 counter$count = 65641;
	#10 counter$count = 65642;
	#10 counter$count = 65643;
	#10 counter$count = 65644;
	#10 counter$count = 65645;
	#10 counter$count = 65646;
	#10 counter$count = 65647;
	#10 counter$count = 65648;
	#10 counter$count = 65649;
	#10 counter$count = 65650;
	#10 counter$count = 65651;
	#10 counter$count = 65652;
	#10 counter$count = 65653;
	#10 counter$count = 65654;
	#10 counter$count = 65655;
	#10 counter$count = 65656;
	#10 counter$count = 65657;
	#10 counter$count = 65658;
	#10 counter$count = 65659;
	#10 counter$count = 65660;
	#10 counter$count = 65661;
	#10 counter$count = 65662;
	#10 counter$count = 65663;
	#10 counter$count = 65664;
	#10 counter$count = 65665;
	#10 counter$count = 65666;
	#10 counter$count = 65667;
	#10 counter$count = 65668;
	#10 counter$count = 65669;
	#10 counter$count = 65670;
	#10 counter$count = 65671;
	#10 counter$count = 65672;
	#10 counter$count = 65673;
	#10 counter$count = 65674;
	#10 counter$count = 65675;
	#10 counter$count = 65676;
	#10 counter$count = 65677;
	#10 counter$count = 65678;
	#10 counter$count = 65679;
	#10 counter$count = 65680;
	#10 counter$count = 65681;
	#10 counter$count = 65682;
	#10 counter$count = 65683;
	#10 counter$count = 65684;
	#10 counter$count = 65685;
	#10 counter$count = 65686;
	#10 counter$count = 65687;
	#10 counter$count = 65688;
	#10 counter$count = 65689;
	#10 counter$count = 65690;
	#10 counter$count = 65691;
	#10 counter$count = 65692;
	#10 counter$count = 65693;
	#10 counter$count = 65694;
	#10 counter$count = 65695;
	#10 counter$count = 65696;
	#10 counter$count = 65697;
	#10 counter$count = 65698;
	#10 counter$count = 65699;
	#10 counter$count = 65700;
	#10 counter$count = 65701;
	#10 counter$count = 65702;
	#10 counter$count = 65703;
	#10 counter$count = 65704;
	#10 counter$count = 65705;
	#10 counter$count = 65706;
	#10 counter$count = 65707;
	#10 counter$count = 65708;
	#10 counter$count = 65709;
	#10 counter$count = 65710;
	#10 counter$count = 65711;
	#10 counter$count = 65712;
	#10 counter$count = 65713;
	#10 counter$count = 65714;
	#10 counter$count = 65715;
	#10 counter$count = 65716;
	#10 counter$count = 65717;
	#10 counter$count = 65718;
	#10 counter$count = 65719;
	#10 counter$count = 65720;
	#10 counter$count = 65721;
	#10 counter$count = 65722;
	#10 counter$count = 65723;
	#10 counter$count = 65724;
	#10 counter$count = 65725;
	#10 counter$count = 65726;
	#10 counter$count = 65727;
	#10 counter$count = 65728;
	#10 counter$count = 65729;
	#10 counter$count = 65730;
	#10 counter$count = 65731;
	#10 counter$count = 65732;
	#10 counter$count = 65733;
	#10 counter$count = 65734;
	#10 counter$count = 65735;
	#10 counter$count = 65736;
	#10 counter$count = 65737;
	#10 counter$count = 65738;
	#10 counter$count = 65739;
	#10 counter$count = 65740;
	#10 counter$count = 65741;
	#10 counter$count = 65742;
	#10 counter$count = 65743;
	#10 counter$count = 65744;
	#10 counter$count = 65745;
	#10 counter$count = 65746;
	#10 counter$count = 65747;
	#10 counter$count = 65748;
	#10 counter$count = 65749;
	#10 counter$count = 65750;
	#10 counter$count = 65751;
	#10 counter$count = 65752;
	#10 counter$count = 65753;
	#10 counter$count = 65754;
	#10 counter$count = 65755;
	#10 counter$count = 65756;
	#10 counter$count = 65757;
	#10 counter$count = 65758;
	#10 counter$count = 65759;
	#10 counter$count = 65760;
	#10 counter$count = 65761;
	#10 counter$count = 65762;
	#10 counter$count = 65763;
	#10 counter$count = 65764;
	#10 counter$count = 65765;
	#10 counter$count = 65766;
	#10 counter$count = 65767;
	#10 counter$count = 65768;
	#10 counter$count = 65769;
	#10 counter$count = 65770;
	#10 counter$count = 65771;
	#10 counter$count = 65772;
	#10 counter$count = 65773;
	#10 counter$count = 65774;
	#10 counter$count = 65775;
	#10 counter$count = 65776;
	#10 counter$count = 65777;
	#10 counter$count = 65778;
	#10 counter$count = 65779;
	#10 counter$count = 65780;
	#10 counter$count = 65781;
	#10 counter$count = 65782;
	#10 counter$count = 65783;
	#10 counter$count = 65784;
	#10 counter$count = 65785;
	#10 counter$count = 65786;
	#10 counter$count = 65787;
	#10 counter$count = 65788;
	#10 counter$count = 65789;
	#10 counter$count = 65790;
	#10 counter$count = 65791;
	#10 counter$count = 65792;
	#10 counter$count = 65793;
	#10 counter$count = 65794;
	#10 counter$count = 65795;
	#10 counter$count = 65796;
	#10 counter$count = 65797;
	#10 counter$count = 65798;
	#10 counter$count = 65799;
	#10 counter$count = 65800;
	#10 counter$count = 65801;
	#10 counter$count = 65802;
	#10 counter$count = 65803;
	#10 counter$count = 65804;
	#10 counter$count = 65805;
	#10 counter$count = 65806;
	#10 counter$count = 65807;
	#10 counter$count = 65808;
	#10 counter$count = 65809;
	#10 counter$count = 65810;
	#10 counter$count = 65811;
	#10 counter$count = 65812;
	#10 counter$count = 65813;
	#10 counter$count = 65814;
	#10 counter$count = 65815;
	#10 counter$count = 65816;
	#10 counter$count = 65817;
	#10 counter$count = 65818;
	#10 counter$count = 65819;
	#10 counter$count = 65820;
	#10 counter$count = 65821;
	#10 counter$count = 65822;
	#10 counter$count = 65823;
	#10 counter$count = 65824;
	#10 counter$count = 65825;
	#10 counter$count = 65826;
	#10 counter$count = 65827;
	#10 counter$count = 65828;
	#10 counter$count = 65829;
	#10 counter$count = 65830;
	#10 counter$count = 65831;
	#10 counter$count = 65832;
	#10 counter$count = 65833;
	#10 counter$count = 65834;
	#10 counter$count = 65835;
	#10 counter$count = 65836;
	#10 counter$count = 65837;
	#10 counter$count = 65838;
	#10 counter$count = 65839;
	#10 counter$count = 65840;
	#10 counter$count = 65841;
	#10 counter$count = 65842;
	#10 counter$count = 65843;
	#10 counter$count = 65844;
	#10 counter$count = 65845;
	#10 counter$count = 65846;
	#10 counter$count = 65847;
	#10 counter$count = 65848;
	#10 counter$count = 65849;
	#10 counter$count = 65850;
	#10 counter$count = 65851;
	#10 counter$count = 65852;
	#10 counter$count = 65853;
	#10 counter$count = 65854;
	#10 counter$count = 65855;
	#10 counter$count = 65856;
	#10 counter$count = 65857;
	#10 counter$count = 65858;
	#10 counter$count = 65859;
	#10 counter$count = 65860;
	#10 counter$count = 65861;
	#10 counter$count = 65862;
	#10 counter$count = 65863;
	#10 counter$count = 65864;
	#10 counter$count = 65865;
	#10 counter$count = 65866;
	#10 counter$count = 65867;
	#10 counter$count = 65868;
	#10 counter$count = 65869;
	#10 counter$count = 65870;
	#10 counter$count = 65871;
	#10 counter$count = 65872;
	#10 counter$count = 65873;
	#10 counter$count = 65874;
	#10 counter$count = 65875;
	#10 counter$count = 65876;
	#10 counter$count = 65877;
	#10 counter$count = 65878;
	#10 counter$count = 65879;
	#10 counter$count = 65880;
	#10 counter$count = 65881;
	#10 counter$count = 65882;
	#10 counter$count = 65883;
	#10 counter$count = 65884;
	#10 counter$count = 65885;
	#10 counter$count = 65886;
	#10 counter$count = 65887;
	#10 counter$count = 65888;
	#10 counter$count = 65889;
	#10 counter$count = 65890;
	#10 counter$count = 65891;
	#10 counter$count = 65892;
	#10 counter$count = 65893;
	#10 counter$count = 65894;
	#10 counter$count = 65895;
	#10 counter$count = 65896;
	#10 counter$count = 65897;
	#10 counter$count = 65898;
	#10 counter$count = 65899;
	#10 counter$count = 65900;
	#10 counter$count = 65901;
	#10 counter$count = 65902;
	#10 counter$count = 65903;
	#10 counter$count = 65904;
	#10 counter$count = 65905;
	#10 counter$count = 65906;
	#10 counter$count = 65907;
	#10 counter$count = 65908;
	#10 counter$count = 65909;
	#10 counter$count = 65910;
	#10 counter$count = 65911;
	#10 counter$count = 65912;
	#10 counter$count = 65913;
	#10 counter$count = 65914;
	#10 counter$count = 65915;
	#10 counter$count = 65916;
	#10 counter$count = 65917;
	#10 counter$count = 65918;
	#10 counter$count = 65919;
	#10 counter$count = 65920;
	#10 counter$count = 65921;
	#10 counter$count = 65922;
	#10 counter$count = 65923;
	#10 counter$count = 65924;
	#10 counter$count = 65925;
	#10 counter$count = 65926;
	#10 counter$count = 65927;
	#10 counter$count = 65928;
	#10 counter$count = 65929;
	#10 counter$count = 65930;
	#10 counter$count = 65931;
	#10 counter$count = 65932;
	#10 counter$count = 65933;
	#10 counter$count = 65934;
	#10 counter$count = 65935;
	#10 counter$count = 65936;
	#10 counter$count = 65937;
	#10 counter$count = 65938;
	#10 counter$count = 65939;
	#10 counter$count = 65940;
	#10 counter$count = 65941;
	#10 counter$count = 65942;
	#10 counter$count = 65943;
	#10 counter$count = 65944;
	#10 counter$count = 65945;
	#10 counter$count = 65946;
	#10 counter$count = 65947;
	#10 counter$count = 65948;
	#10 counter$count = 65949;
	#10 counter$count = 65950;
	#10 counter$count = 65951;
	#10 counter$count = 65952;
	#10 counter$count = 65953;
	#10 counter$count = 65954;
	#10 counter$count = 65955;
	#10 counter$count = 65956;
	#10 counter$count = 65957;
	#10 counter$count = 65958;
	#10 counter$count = 65959;
	#10 counter$count = 65960;
	#10 counter$count = 65961;
	#10 counter$count = 65962;
	#10 counter$count = 65963;
	#10 counter$count = 65964;
	#10 counter$count = 65965;
	#10 counter$count = 65966;
	#10 counter$count = 65967;
	#10 counter$count = 65968;
	#10 counter$count = 65969;
	#10 counter$count = 65970;
	#10 counter$count = 65971;
	#10 counter$count = 65972;
	#10 counter$count = 65973;
	#10 counter$count = 65974;
	#10 counter$count = 65975;
	#10 counter$count = 65976;
	#10 counter$count = 65977;
	#10 counter$count = 65978;
	#10 counter$count = 65979;
	#10 counter$count = 65980;
	#10 counter$count = 65981;
	#10 counter$count = 65982;
	#10 counter$count = 65983;
	#10 counter$count = 65984;
	#10 counter$count = 65985;
	#10 counter$count = 65986;
	#10 counter$count = 65987;
	#10 counter$count = 65988;
	#10 counter$count = 65989;
	#10 counter$count = 65990;
	#10 counter$count = 65991;
	#10 counter$count = 65992;
	#10 counter$count = 65993;
	#10 counter$count = 65994;
	#10 counter$count = 65995;
	#10 counter$count = 65996;
	#10 counter$count = 65997;
	#10 counter$count = 65998;
	#10 counter$count = 65999;
	#10 counter$count = 66000;
	#10 counter$count = 66001;
	#10 counter$count = 66002;
	#10 counter$count = 66003;
	#10 counter$count = 66004;
	#10 counter$count = 66005;
	#10 counter$count = 66006;
	#10 counter$count = 66007;
	#10 counter$count = 66008;
	#10 counter$count = 66009;
	#10 counter$count = 66010;
	#10 counter$count = 66011;
	#10 counter$count = 66012;
	#10 counter$count = 66013;
	#10 counter$count = 66014;
	#10 counter$count = 66015;
	#10 counter$count = 66016;
	#10 counter$count = 66017;
	#10 counter$count = 66018;
	#10 counter$count = 66019;
	#10 counter$count = 66020;
	#10 counter$count = 66021;
	#10 counter$count = 66022;
	#10 counter$count = 66023;
	#10 counter$count = 66024;
	#10 counter$count = 66025;
	#10 counter$count = 66026;
	#10 counter$count = 66027;
	#10 counter$count = 66028;
	#10 counter$count = 66029;
	#10 counter$count = 66030;
	#10 counter$count = 66031;
	#10 counter$count = 66032;
	#10 counter$count = 66033;
	#10 counter$count = 66034;
	#10 counter$count = 66035;
	#10 counter$count = 66036;
	#10 counter$count = 66037;
	#10 counter$count = 66038;
	#10 counter$count = 66039;
	#10 counter$count = 66040;
	#10 counter$count = 66041;
	#10 counter$count = 66042;
	#10 counter$count = 66043;
	#10 counter$count = 66044;
	#10 counter$count = 66045;
	#10 counter$count = 66046;
	#10 counter$count = 66047;
	#10 counter$count = 66048;
	#10 counter$count = 66049;
	#10 counter$count = 66050;
	#10 counter$count = 66051;
	#10 counter$count = 66052;
	#10 counter$count = 66053;
	#10 counter$count = 66054;
	#10 counter$count = 66055;
	#10 counter$count = 66056;
	#10 counter$count = 66057;
	#10 counter$count = 66058;
	#10 counter$count = 66059;
	#10 counter$count = 66060;
	#10 counter$count = 66061;
	#10 counter$count = 66062;
	#10 counter$count = 66063;
	#10 counter$count = 66064;
	#10 counter$count = 66065;
	#10 counter$count = 66066;
	#10 counter$count = 66067;
	#10 counter$count = 66068;
	#10 counter$count = 66069;
	#10 counter$count = 66070;
	#10 counter$count = 66071;
	#10 counter$count = 66072;
	#10 counter$count = 66073;
	#10 counter$count = 66074;
	#10 counter$count = 66075;
	#10 counter$count = 66076;
	#10 counter$count = 66077;
	#10 counter$count = 66078;
	#10 counter$count = 66079;
	#10 counter$count = 66080;
	#10 counter$count = 66081;
	#10 counter$count = 66082;
	#10 counter$count = 66083;
	#10 counter$count = 66084;
	#10 counter$count = 66085;
	#10 counter$count = 66086;
	#10 counter$count = 66087;
	#10 counter$count = 66088;
	#10 counter$count = 66089;
	#10 counter$count = 66090;
	#10 counter$count = 66091;
	#10 counter$count = 66092;
	#10 counter$count = 66093;
	#10 counter$count = 66094;
	#10 counter$count = 66095;
	#10 counter$count = 66096;
	#10 counter$count = 66097;
	#10 counter$count = 66098;
	#10 counter$count = 66099;
	#10 counter$count = 66100;
	#10 counter$count = 66101;
	#10 counter$count = 66102;
	#10 counter$count = 66103;
	#10 counter$count = 66104;
	#10 counter$count = 66105;
	#10 counter$count = 66106;
	#10 counter$count = 66107;
	#10 counter$count = 66108;
	#10 counter$count = 66109;
	#10 counter$count = 66110;
	#10 counter$count = 66111;
	#10 counter$count = 66112;
	#10 counter$count = 66113;
	#10 counter$count = 66114;
	#10 counter$count = 66115;
	#10 counter$count = 66116;
	#10 counter$count = 66117;
	#10 counter$count = 66118;
	#10 counter$count = 66119;
	#10 counter$count = 66120;
	#10 counter$count = 66121;
	#10 counter$count = 66122;
	#10 counter$count = 66123;
	#10 counter$count = 66124;
	#10 counter$count = 66125;
	#10 counter$count = 66126;
	#10 counter$count = 66127;
	#10 counter$count = 66128;
	#10 counter$count = 66129;
	#10 counter$count = 66130;
	#10 counter$count = 66131;
	#10 counter$count = 66132;
	#10 counter$count = 66133;
	#10 counter$count = 66134;
	#10 counter$count = 66135;
	#10 counter$count = 66136;
	#10 counter$count = 66137;
	#10 counter$count = 66138;
	#10 counter$count = 66139;
	#10 counter$count = 66140;
	#10 counter$count = 66141;
	#10 counter$count = 66142;
	#10 counter$count = 66143;
	#10 counter$count = 66144;
	#10 counter$count = 66145;
	#10 counter$count = 66146;
	#10 counter$count = 66147;
	#10 counter$count = 66148;
	#10 counter$count = 66149;
	#10 counter$count = 66150;
	#10 counter$count = 66151;
	#10 counter$count = 66152;
	#10 counter$count = 66153;
	#10 counter$count = 66154;
	#10 counter$count = 66155;
	#10 counter$count = 66156;
	#10 counter$count = 66157;
	#10 counter$count = 66158;
	#10 counter$count = 66159;
	#10 counter$count = 66160;
	#10 counter$count = 66161;
	#10 counter$count = 66162;
	#10 counter$count = 66163;
	#10 counter$count = 66164;
	#10 counter$count = 66165;
	#10 counter$count = 66166;
	#10 counter$count = 66167;
	#10 counter$count = 66168;
	#10 counter$count = 66169;
	#10 counter$count = 66170;
	#10 counter$count = 66171;
	#10 counter$count = 66172;
	#10 counter$count = 66173;
	#10 counter$count = 66174;
	#10 counter$count = 66175;
	#10 counter$count = 66176;
	#10 counter$count = 66177;
	#10 counter$count = 66178;
	#10 counter$count = 66179;
	#10 counter$count = 66180;
	#10 counter$count = 66181;
	#10 counter$count = 66182;
	#10 counter$count = 66183;
	#10 counter$count = 66184;
	#10 counter$count = 66185;
	#10 counter$count = 66186;
	#10 counter$count = 66187;
	#10 counter$count = 66188;
	#10 counter$count = 66189;
	#10 counter$count = 66190;
	#10 counter$count = 66191;
	#10 counter$count = 66192;
	#10 counter$count = 66193;
	#10 counter$count = 66194;
	#10 counter$count = 66195;
	#10 counter$count = 66196;
	#10 counter$count = 66197;
	#10 counter$count = 66198;
	#10 counter$count = 66199;
	#10 counter$count = 66200;
	#10 counter$count = 66201;
	#10 counter$count = 66202;
	#10 counter$count = 66203;
	#10 counter$count = 66204;
	#10 counter$count = 66205;
	#10 counter$count = 66206;
	#10 counter$count = 66207;
	#10 counter$count = 66208;
	#10 counter$count = 66209;
	#10 counter$count = 66210;
	#10 counter$count = 66211;
	#10 counter$count = 66212;
	#10 counter$count = 66213;
	#10 counter$count = 66214;
	#10 counter$count = 66215;
	#10 counter$count = 66216;
	#10 counter$count = 66217;
	#10 counter$count = 66218;
	#10 counter$count = 66219;
	#10 counter$count = 66220;
	#10 counter$count = 66221;
	#10 counter$count = 66222;
	#10 counter$count = 66223;
	#10 counter$count = 66224;
	#10 counter$count = 66225;
	#10 counter$count = 66226;
	#10 counter$count = 66227;
	#10 counter$count = 66228;
	#10 counter$count = 66229;
	#10 counter$count = 66230;
	#10 counter$count = 66231;
	#10 counter$count = 66232;
	#10 counter$count = 66233;
	#10 counter$count = 66234;
	#10 counter$count = 66235;
	#10 counter$count = 66236;
	#10 counter$count = 66237;
	#10 counter$count = 66238;
	#10 counter$count = 66239;
	#10 counter$count = 66240;
	#10 counter$count = 66241;
	#10 counter$count = 66242;
	#10 counter$count = 66243;
	#10 counter$count = 66244;
	#10 counter$count = 66245;
	#10 counter$count = 66246;
	#10 counter$count = 66247;
	#10 counter$count = 66248;
	#10 counter$count = 66249;
	#10 counter$count = 66250;
	#10 counter$count = 66251;
	#10 counter$count = 66252;
	#10 counter$count = 66253;
	#10 counter$count = 66254;
	#10 counter$count = 66255;
	#10 counter$count = 66256;
	#10 counter$count = 66257;
	#10 counter$count = 66258;
	#10 counter$count = 66259;
	#10 counter$count = 66260;
	#10 counter$count = 66261;
	#10 counter$count = 66262;
	#10 counter$count = 66263;
	#10 counter$count = 66264;
	#10 counter$count = 66265;
	#10 counter$count = 66266;
	#10 counter$count = 66267;
	#10 counter$count = 66268;
	#10 counter$count = 66269;
	#10 counter$count = 66270;
	#10 counter$count = 66271;
	#10 counter$count = 66272;
	#10 counter$count = 66273;
	#10 counter$count = 66274;
	#10 counter$count = 66275;
	#10 counter$count = 66276;
	#10 counter$count = 66277;
	#10 counter$count = 66278;
	#10 counter$count = 66279;
	#10 counter$count = 66280;
	#10 counter$count = 66281;
	#10 counter$count = 66282;
	#10 counter$count = 66283;
	#10 counter$count = 66284;
	#10 counter$count = 66285;
	#10 counter$count = 66286;
	#10 counter$count = 66287;
	#10 counter$count = 66288;
	#10 counter$count = 66289;
	#10 counter$count = 66290;
	#10 counter$count = 66291;
	#10 counter$count = 66292;
	#10 counter$count = 66293;
	#10 counter$count = 66294;
	#10 counter$count = 66295;
	#10 counter$count = 66296;
	#10 counter$count = 66297;
	#10 counter$count = 66298;
	#10 counter$count = 66299;
	#10 counter$count = 66300;
	#10 counter$count = 66301;
	#10 counter$count = 66302;
	#10 counter$count = 66303;
	#10 counter$count = 66304;
	#10 counter$count = 66305;
	#10 counter$count = 66306;
	#10 counter$count = 66307;
	#10 counter$count = 66308;
	#10 counter$count = 66309;
	#10 counter$count = 66310;
	#10 counter$count = 66311;
	#10 counter$count = 66312;
	#10 counter$count = 66313;
	#10 counter$count = 66314;
	#10 counter$count = 66315;
	#10 counter$count = 66316;
	#10 counter$count = 66317;
	#10 counter$count = 66318;
	#10 counter$count = 66319;
	#10 counter$count = 66320;
	#10 counter$count = 66321;
	#10 counter$count = 66322;
	#10 counter$count = 66323;
	#10 counter$count = 66324;
	#10 counter$count = 66325;
	#10 counter$count = 66326;
	#10 counter$count = 66327;
	#10 counter$count = 66328;
	#10 counter$count = 66329;
	#10 counter$count = 66330;
	#10 counter$count = 66331;
	#10 counter$count = 66332;
	#10 counter$count = 66333;
	#10 counter$count = 66334;
	#10 counter$count = 66335;
	#10 counter$count = 66336;
	#10 counter$count = 66337;
	#10 counter$count = 66338;
	#10 counter$count = 66339;
	#10 counter$count = 66340;
	#10 counter$count = 66341;
	#10 counter$count = 66342;
	#10 counter$count = 66343;
	#10 counter$count = 66344;
	#10 counter$count = 66345;
	#10 counter$count = 66346;
	#10 counter$count = 66347;
	#10 counter$count = 66348;
	#10 counter$count = 66349;
	#10 counter$count = 66350;
	#10 counter$count = 66351;
	#10 counter$count = 66352;
	#10 counter$count = 66353;
	#10 counter$count = 66354;
	#10 counter$count = 66355;
	#10 counter$count = 66356;
	#10 counter$count = 66357;
	#10 counter$count = 66358;
	#10 counter$count = 66359;
	#10 counter$count = 66360;
	#10 counter$count = 66361;
	#10 counter$count = 66362;
	#10 counter$count = 66363;
	#10 counter$count = 66364;
	#10 counter$count = 66365;
	#10 counter$count = 66366;
	#10 counter$count = 66367;
	#10 counter$count = 66368;
	#10 counter$count = 66369;
	#10 counter$count = 66370;
	#10 counter$count = 66371;
	#10 counter$count = 66372;
	#10 counter$count = 66373;
	#10 counter$count = 66374;
	#10 counter$count = 66375;
	#10 counter$count = 66376;
	#10 counter$count = 66377;
	#10 counter$count = 66378;
	#10 counter$count = 66379;
	#10 counter$count = 66380;
	#10 counter$count = 66381;
	#10 counter$count = 66382;
	#10 counter$count = 66383;
	#10 counter$count = 66384;
	#10 counter$count = 66385;
	#10 counter$count = 66386;
	#10 counter$count = 66387;
	#10 counter$count = 66388;
	#10 counter$count = 66389;
	#10 counter$count = 66390;
	#10 counter$count = 66391;
	#10 counter$count = 66392;
	#10 counter$count = 66393;
	#10 counter$count = 66394;
	#10 counter$count = 66395;
	#10 counter$count = 66396;
	#10 counter$count = 66397;
	#10 counter$count = 66398;
	#10 counter$count = 66399;
	#10 counter$count = 66400;
	#10 counter$count = 66401;
	#10 counter$count = 66402;
	#10 counter$count = 66403;
	#10 counter$count = 66404;
	#10 counter$count = 66405;
	#10 counter$count = 66406;
	#10 counter$count = 66407;
	#10 counter$count = 66408;
	#10 counter$count = 66409;
	#10 counter$count = 66410;
	#10 counter$count = 66411;
	#10 counter$count = 66412;
	#10 counter$count = 66413;
	#10 counter$count = 66414;
	#10 counter$count = 66415;
	#10 counter$count = 66416;
	#10 counter$count = 66417;
	#10 counter$count = 66418;
	#10 counter$count = 66419;
	#10 counter$count = 66420;
	#10 counter$count = 66421;
	#10 counter$count = 66422;
	#10 counter$count = 66423;
	#10 counter$count = 66424;
	#10 counter$count = 66425;
	#10 counter$count = 66426;
	#10 counter$count = 66427;
	#10 counter$count = 66428;
	#10 counter$count = 66429;
	#10 counter$count = 66430;
	#10 counter$count = 66431;
	#10 counter$count = 66432;
	#10 counter$count = 66433;
	#10 counter$count = 66434;
	#10 counter$count = 66435;
	#10 counter$count = 66436;
	#10 counter$count = 66437;
	#10 counter$count = 66438;
	#10 counter$count = 66439;
	#10 counter$count = 66440;
	#10 counter$count = 66441;
	#10 counter$count = 66442;
	#10 counter$count = 66443;
	#10 counter$count = 66444;
	#10 counter$count = 66445;
	#10 counter$count = 66446;
	#10 counter$count = 66447;
	#10 counter$count = 66448;
	#10 counter$count = 66449;
	#10 counter$count = 66450;
	#10 counter$count = 66451;
	#10 counter$count = 66452;
	#10 counter$count = 66453;
	#10 counter$count = 66454;
	#10 counter$count = 66455;
	#10 counter$count = 66456;
	#10 counter$count = 66457;
	#10 counter$count = 66458;
	#10 counter$count = 66459;
	#10 counter$count = 66460;
	#10 counter$count = 66461;
	#10 counter$count = 66462;
	#10 counter$count = 66463;
	#10 counter$count = 66464;
	#10 counter$count = 66465;
	#10 counter$count = 66466;
	#10 counter$count = 66467;
	#10 counter$count = 66468;
	#10 counter$count = 66469;
	#10 counter$count = 66470;
	#10 counter$count = 66471;
	#10 counter$count = 66472;
	#10 counter$count = 66473;
	#10 counter$count = 66474;
	#10 counter$count = 66475;
	#10 counter$count = 66476;
	#10 counter$count = 66477;
	#10 counter$count = 66478;
	#10 counter$count = 66479;
	#10 counter$count = 66480;
	#10 counter$count = 66481;
	#10 counter$count = 66482;
	#10 counter$count = 66483;
	#10 counter$count = 66484;
	#10 counter$count = 66485;
	#10 counter$count = 66486;
	#10 counter$count = 66487;
	#10 counter$count = 66488;
	#10 counter$count = 66489;
	#10 counter$count = 66490;
	#10 counter$count = 66491;
	#10 counter$count = 66492;
	#10 counter$count = 66493;
	#10 counter$count = 66494;
	#10 counter$count = 66495;
	#10 counter$count = 66496;
	#10 counter$count = 66497;
	#10 counter$count = 66498;
	#10 counter$count = 66499;
	#10 counter$count = 66500;
	#10 counter$count = 66501;
	#10 counter$count = 66502;
	#10 counter$count = 66503;
	#10 counter$count = 66504;
	#10 counter$count = 66505;
	#10 counter$count = 66506;
	#10 counter$count = 66507;
	#10 counter$count = 66508;
	#10 counter$count = 66509;
	#10 counter$count = 66510;
	#10 counter$count = 66511;
	#10 counter$count = 66512;
	#10 counter$count = 66513;
	#10 counter$count = 66514;
	#10 counter$count = 66515;
	#10 counter$count = 66516;
	#10 counter$count = 66517;
	#10 counter$count = 66518;
	#10 counter$count = 66519;
	#10 counter$count = 66520;
	#10 counter$count = 66521;
	#10 counter$count = 66522;
	#10 counter$count = 66523;
	#10 counter$count = 66524;
	#10 counter$count = 66525;
	#10 counter$count = 66526;
	#10 counter$count = 66527;
	#10 counter$count = 66528;
	#10 counter$count = 66529;
	#10 counter$count = 66530;
	#10 counter$count = 66531;
	#10 counter$count = 66532;
	#10 counter$count = 66533;
	#10 counter$count = 66534;
	#10 counter$count = 66535;
	#10 counter$count = 66536;
	#10 counter$count = 66537;
	#10 counter$count = 66538;
	#10 counter$count = 66539;
	#10 counter$count = 66540;
	#10 counter$count = 66541;
	#10 counter$count = 66542;
	#10 counter$count = 66543;
	#10 counter$count = 66544;
	#10 counter$count = 66545;
	#10 counter$count = 66546;
	#10 counter$count = 66547;
	#10 counter$count = 66548;
	#10 counter$count = 66549;
	#10 counter$count = 66550;
	#10 counter$count = 66551;
	#10 counter$count = 66552;
	#10 counter$count = 66553;
	#10 counter$count = 66554;
	#10 counter$count = 66555;
	#10 counter$count = 66556;
	#10 counter$count = 66557;
	#10 counter$count = 66558;
	#10 counter$count = 66559;
	#10 counter$count = 66560;
	#10 counter$count = 66561;
	#10 counter$count = 66562;
	#10 counter$count = 66563;
	#10 counter$count = 66564;
	#10 counter$count = 66565;
	#10 counter$count = 66566;
	#10 counter$count = 66567;
	#10 counter$count = 66568;
	#10 counter$count = 66569;
	#10 counter$count = 66570;
	#10 counter$count = 66571;
	#10 counter$count = 66572;
	#10 counter$count = 66573;
	#10 counter$count = 66574;
	#10 counter$count = 66575;
	#10 counter$count = 66576;
	#10 counter$count = 66577;
	#10 counter$count = 66578;
	#10 counter$count = 66579;
	#10 counter$count = 66580;
	#10 counter$count = 66581;
	#10 counter$count = 66582;
	#10 counter$count = 66583;
	#10 counter$count = 66584;
	#10 counter$count = 66585;
	#10 counter$count = 66586;
	#10 counter$count = 66587;
	#10 counter$count = 66588;
	#10 counter$count = 66589;
	#10 counter$count = 66590;
	#10 counter$count = 66591;
	#10 counter$count = 66592;
	#10 counter$count = 66593;
	#10 counter$count = 66594;
	#10 counter$count = 66595;
	#10 counter$count = 66596;
	#10 counter$count = 66597;
	#10 counter$count = 66598;
	#10 counter$count = 66599;
	#10 counter$count = 66600;
	#10 counter$count = 66601;
	#10 counter$count = 66602;
	#10 counter$count = 66603;
	#10 counter$count = 66604;
	#10 counter$count = 66605;
	#10 counter$count = 66606;
	#10 counter$count = 66607;
	#10 counter$count = 66608;
	#10 counter$count = 66609;
	#10 counter$count = 66610;
	#10 counter$count = 66611;
	#10 counter$count = 66612;
	#10 counter$count = 66613;
	#10 counter$count = 66614;
	#10 counter$count = 66615;
	#10 counter$count = 66616;
	#10 counter$count = 66617;
	#10 counter$count = 66618;
	#10 counter$count = 66619;
	#10 counter$count = 66620;
	#10 counter$count = 66621;
	#10 counter$count = 66622;
	#10 counter$count = 66623;
	#10 counter$count = 66624;
	#10 counter$count = 66625;
	#10 counter$count = 66626;
	#10 counter$count = 66627;
	#10 counter$count = 66628;
	#10 counter$count = 66629;
	#10 counter$count = 66630;
	#10 counter$count = 66631;
	#10 counter$count = 66632;
	#10 counter$count = 66633;
	#10 counter$count = 66634;
	#10 counter$count = 66635;
	#10 counter$count = 66636;
	#10 counter$count = 66637;
	#10 counter$count = 66638;
	#10 counter$count = 66639;
	#10 counter$count = 66640;
	#10 counter$count = 66641;
	#10 counter$count = 66642;
	#10 counter$count = 66643;
	#10 counter$count = 66644;
	#10 counter$count = 66645;
	#10 counter$count = 66646;
	#10 counter$count = 66647;
	#10 counter$count = 66648;
	#10 counter$count = 66649;
	#10 counter$count = 66650;
	#10 counter$count = 66651;
	#10 counter$count = 66652;
	#10 counter$count = 66653;
	#10 counter$count = 66654;
	#10 counter$count = 66655;
	#10 counter$count = 66656;
	#10 counter$count = 66657;
	#10 counter$count = 66658;
	#10 counter$count = 66659;
	#10 counter$count = 66660;
	#10 counter$count = 66661;
	#10 counter$count = 66662;
	#10 counter$count = 66663;
	#10 counter$count = 66664;
	#10 counter$count = 66665;
	#10 counter$count = 66666;
	#10 counter$count = 66667;
	#10 counter$count = 66668;
	#10 counter$count = 66669;
	#10 counter$count = 66670;
	#10 counter$count = 66671;
	#10 counter$count = 66672;
	#10 counter$count = 66673;
	#10 counter$count = 66674;
	#10 counter$count = 66675;
	#10 counter$count = 66676;
	#10 counter$count = 66677;
	#10 counter$count = 66678;
	#10 counter$count = 66679;
	#10 counter$count = 66680;
	#10 counter$count = 66681;
	#10 counter$count = 66682;
	#10 counter$count = 66683;
	#10 counter$count = 66684;
	#10 counter$count = 66685;
	#10 counter$count = 66686;
	#10 counter$count = 66687;
	#10 counter$count = 66688;
	#10 counter$count = 66689;
	#10 counter$count = 66690;
	#10 counter$count = 66691;
	#10 counter$count = 66692;
	#10 counter$count = 66693;
	#10 counter$count = 66694;
	#10 counter$count = 66695;
	#10 counter$count = 66696;
	#10 counter$count = 66697;
	#10 counter$count = 66698;
	#10 counter$count = 66699;
	#10 counter$count = 66700;
	#10 counter$count = 66701;
	#10 counter$count = 66702;
	#10 counter$count = 66703;
	#10 counter$count = 66704;
	#10 counter$count = 66705;
	#10 counter$count = 66706;
	#10 counter$count = 66707;
	#10 counter$count = 66708;
	#10 counter$count = 66709;
	#10 counter$count = 66710;
	#10 counter$count = 66711;
	#10 counter$count = 66712;
	#10 counter$count = 66713;
	#10 counter$count = 66714;
	#10 counter$count = 66715;
	#10 counter$count = 66716;
	#10 counter$count = 66717;
	#10 counter$count = 66718;
	#10 counter$count = 66719;
	#10 counter$count = 66720;
	#10 counter$count = 66721;
	#10 counter$count = 66722;
	#10 counter$count = 66723;
	#10 counter$count = 66724;
	#10 counter$count = 66725;
	#10 counter$count = 66726;
	#10 counter$count = 66727;
	#10 counter$count = 66728;
	#10 counter$count = 66729;
	#10 counter$count = 66730;
	#10 counter$count = 66731;
	#10 counter$count = 66732;
	#10 counter$count = 66733;
	#10 counter$count = 66734;
	#10 counter$count = 66735;
	#10 counter$count = 66736;
	#10 counter$count = 66737;
	#10 counter$count = 66738;
	#10 counter$count = 66739;
	#10 counter$count = 66740;
	#10 counter$count = 66741;
	#10 counter$count = 66742;
	#10 counter$count = 66743;
	#10 counter$count = 66744;
	#10 counter$count = 66745;
	#10 counter$count = 66746;
	#10 counter$count = 66747;
	#10 counter$count = 66748;
	#10 counter$count = 66749;
	#10 counter$count = 66750;
	#10 counter$count = 66751;
	#10 counter$count = 66752;
	#10 counter$count = 66753;
	#10 counter$count = 66754;
	#10 counter$count = 66755;
	#10 counter$count = 66756;
	#10 counter$count = 66757;
	#10 counter$count = 66758;
	#10 counter$count = 66759;
	#10 counter$count = 66760;
	#10 counter$count = 66761;
	#10 counter$count = 66762;
	#10 counter$count = 66763;
	#10 counter$count = 66764;
	#10 counter$count = 66765;
	#10 counter$count = 66766;
	#10 counter$count = 66767;
	#10 counter$count = 66768;
	#10 counter$count = 66769;
	#10 counter$count = 66770;
	#10 counter$count = 66771;
	#10 counter$count = 66772;
	#10 counter$count = 66773;
	#10 counter$count = 66774;
	#10 counter$count = 66775;
	#10 counter$count = 66776;
	#10 counter$count = 66777;
	#10 counter$count = 66778;
	#10 counter$count = 66779;
	#10 counter$count = 66780;
	#10 counter$count = 66781;
	#10 counter$count = 66782;
	#10 counter$count = 66783;
	#10 counter$count = 66784;
	#10 counter$count = 66785;
	#10 counter$count = 66786;
	#10 counter$count = 66787;
	#10 counter$count = 66788;
	#10 counter$count = 66789;
	#10 counter$count = 66790;
	#10 counter$count = 66791;
	#10 counter$count = 66792;
	#10 counter$count = 66793;
	#10 counter$count = 66794;
	#10 counter$count = 66795;
	#10 counter$count = 66796;
	#10 counter$count = 66797;
	#10 counter$count = 66798;
	#10 counter$count = 66799;
	#10 counter$count = 66800;
	#10 counter$count = 66801;
	#10 counter$count = 66802;
	#10 counter$count = 66803;
	#10 counter$count = 66804;
	#10 counter$count = 66805;
	#10 counter$count = 66806;
	#10 counter$count = 66807;
	#10 counter$count = 66808;
	#10 counter$count = 66809;
	#10 counter$count = 66810;
	#10 counter$count = 66811;
	#10 counter$count = 66812;
	#10 counter$count = 66813;
	#10 counter$count = 66814;
	#10 counter$count = 66815;
	#10 counter$count = 66816;
	#10 counter$count = 66817;
	#10 counter$count = 66818;
	#10 counter$count = 66819;
	#10 counter$count = 66820;
	#10 counter$count = 66821;
	#10 counter$count = 66822;
	#10 counter$count = 66823;
	#10 counter$count = 66824;
	#10 counter$count = 66825;
	#10 counter$count = 66826;
	#10 counter$count = 66827;
	#10 counter$count = 66828;
	#10 counter$count = 66829;
	#10 counter$count = 66830;
	#10 counter$count = 66831;
	#10 counter$count = 66832;
	#10 counter$count = 66833;
	#10 counter$count = 66834;
	#10 counter$count = 66835;
	#10 counter$count = 66836;
	#10 counter$count = 66837;
	#10 counter$count = 66838;
	#10 counter$count = 66839;
	#10 counter$count = 66840;
	#10 counter$count = 66841;
	#10 counter$count = 66842;
	#10 counter$count = 66843;
	#10 counter$count = 66844;
	#10 counter$count = 66845;
	#10 counter$count = 66846;
	#10 counter$count = 66847;
	#10 counter$count = 66848;
	#10 counter$count = 66849;
	#10 counter$count = 66850;
	#10 counter$count = 66851;
	#10 counter$count = 66852;
	#10 counter$count = 66853;
	#10 counter$count = 66854;
	#10 counter$count = 66855;
	#10 counter$count = 66856;
	#10 counter$count = 66857;
	#10 counter$count = 66858;
	#10 counter$count = 66859;
	#10 counter$count = 66860;
	#10 counter$count = 66861;
	#10 counter$count = 66862;
	#10 counter$count = 66863;
	#10 counter$count = 66864;
	#10 counter$count = 66865;
	#10 counter$count = 66866;
	#10 counter$count = 66867;
	#10 counter$count = 66868;
	#10 counter$count = 66869;
	#10 counter$count = 66870;
	#10 counter$count = 66871;
	#10 counter$count = 66872;
	#10 counter$count = 66873;
	#10 counter$count = 66874;
	#10 counter$count = 66875;
	#10 counter$count = 66876;
	#10 counter$count = 66877;
	#10 counter$count = 66878;
	#10 counter$count = 66879;
	#10 counter$count = 66880;
	#10 counter$count = 66881;
	#10 counter$count = 66882;
	#10 counter$count = 66883;
	#10 counter$count = 66884;
	#10 counter$count = 66885;
	#10 counter$count = 66886;
	#10 counter$count = 66887;
	#10 counter$count = 66888;
	#10 counter$count = 66889;
	#10 counter$count = 66890;
	#10 counter$count = 66891;
	#10 counter$count = 66892;
	#10 counter$count = 66893;
	#10 counter$count = 66894;
	#10 counter$count = 66895;
	#10 counter$count = 66896;
	#10 counter$count = 66897;
	#10 counter$count = 66898;
	#10 counter$count = 66899;
	#10 counter$count = 66900;
	#10 counter$count = 66901;
	#10 counter$count = 66902;
	#10 counter$count = 66903;
	#10 counter$count = 66904;
	#10 counter$count = 66905;
	#10 counter$count = 66906;
	#10 counter$count = 66907;
	#10 counter$count = 66908;
	#10 counter$count = 66909;
	#10 counter$count = 66910;
	#10 counter$count = 66911;
	#10 counter$count = 66912;
	#10 counter$count = 66913;
	#10 counter$count = 66914;
	#10 counter$count = 66915;
	#10 counter$count = 66916;
	#10 counter$count = 66917;
	#10 counter$count = 66918;
	#10 counter$count = 66919;
	#10 counter$count = 66920;
	#10 counter$count = 66921;
	#10 counter$count = 66922;
	#10 counter$count = 66923;
	#10 counter$count = 66924;
	#10 counter$count = 66925;
	#10 counter$count = 66926;
	#10 counter$count = 66927;
	#10 counter$count = 66928;
	#10 counter$count = 66929;
	#10 counter$count = 66930;
	#10 counter$count = 66931;
	#10 counter$count = 66932;
	#10 counter$count = 66933;
	#10 counter$count = 66934;
	#10 counter$count = 66935;
	#10 counter$count = 66936;
	#10 counter$count = 66937;
	#10 counter$count = 66938;
	#10 counter$count = 66939;
	#10 counter$count = 66940;
	#10 counter$count = 66941;
	#10 counter$count = 66942;
	#10 counter$count = 66943;
	#10 counter$count = 66944;
	#10 counter$count = 66945;
	#10 counter$count = 66946;
	#10 counter$count = 66947;
	#10 counter$count = 66948;
	#10 counter$count = 66949;
	#10 counter$count = 66950;
	#10 counter$count = 66951;
	#10 counter$count = 66952;
	#10 counter$count = 66953;
	#10 counter$count = 66954;
	#10 counter$count = 66955;
	#10 counter$count = 66956;
	#10 counter$count = 66957;
	#10 counter$count = 66958;
	#10 counter$count = 66959;
	#10 counter$count = 66960;
	#10 counter$count = 66961;
	#10 counter$count = 66962;
	#10 counter$count = 66963;
	#10 counter$count = 66964;
	#10 counter$count = 66965;
	#10 counter$count = 66966;
	#10 counter$count = 66967;
	#10 counter$count = 66968;
	#10 counter$count = 66969;
	#10 counter$count = 66970;
	#10 counter$count = 66971;
	#10 counter$count = 66972;
	#10 counter$count = 66973;
	#10 counter$count = 66974;
	#10 counter$count = 66975;
	#10 counter$count = 66976;
	#10 counter$count = 66977;
	#10 counter$count = 66978;
	#10 counter$count = 66979;
	#10 counter$count = 66980;
	#10 counter$count = 66981;
	#10 counter$count = 66982;
	#10 counter$count = 66983;
	#10 counter$count = 66984;
	#10 counter$count = 66985;
	#10 counter$count = 66986;
	#10 counter$count = 66987;
	#10 counter$count = 66988;
	#10 counter$count = 66989;
	#10 counter$count = 66990;
	#10 counter$count = 66991;
	#10 counter$count = 66992;
	#10 counter$count = 66993;
	#10 counter$count = 66994;
	#10 counter$count = 66995;
	#10 counter$count = 66996;
	#10 counter$count = 66997;
	#10 counter$count = 66998;
	#10 counter$count = 66999;
	#10 counter$count = 67000;
	#10 counter$count = 67001;
	#10 counter$count = 67002;
	#10 counter$count = 67003;
	#10 counter$count = 67004;
	#10 counter$count = 67005;
	#10 counter$count = 67006;
	#10 counter$count = 67007;
	#10 counter$count = 67008;
	#10 counter$count = 67009;
	#10 counter$count = 67010;
	#10 counter$count = 67011;
	#10 counter$count = 67012;
	#10 counter$count = 67013;
	#10 counter$count = 67014;
	#10 counter$count = 67015;
	#10 counter$count = 67016;
	#10 counter$count = 67017;
	#10 counter$count = 67018;
	#10 counter$count = 67019;
	#10 counter$count = 67020;
	#10 counter$count = 67021;
	#10 counter$count = 67022;
	#10 counter$count = 67023;
	#10 counter$count = 67024;
	#10 counter$count = 67025;
	#10 counter$count = 67026;
	#10 counter$count = 67027;
	#10 counter$count = 67028;
	#10 counter$count = 67029;
	#10 counter$count = 67030;
	#10 counter$count = 67031;
	#10 counter$count = 67032;
	#10 counter$count = 67033;
	#10 counter$count = 67034;
	#10 counter$count = 67035;
	#10 counter$count = 67036;
	#10 counter$count = 67037;
	#10 counter$count = 67038;
	#10 counter$count = 67039;
	#10 counter$count = 67040;
	#10 counter$count = 67041;
	#10 counter$count = 67042;
	#10 counter$count = 67043;
	#10 counter$count = 67044;
	#10 counter$count = 67045;
	#10 counter$count = 67046;
	#10 counter$count = 67047;
	#10 counter$count = 67048;
	#10 counter$count = 67049;
	#10 counter$count = 67050;
	#10 counter$count = 67051;
	#10 counter$count = 67052;
	#10 counter$count = 67053;
	#10 counter$count = 67054;
	#10 counter$count = 67055;
	#10 counter$count = 67056;
	#10 counter$count = 67057;
	#10 counter$count = 67058;
	#10 counter$count = 67059;
	#10 counter$count = 67060;
	#10 counter$count = 67061;
	#10 counter$count = 67062;
	#10 counter$count = 67063;
	#10 counter$count = 67064;
	#10 counter$count = 67065;
	#10 counter$count = 67066;
	#10 counter$count = 67067;
	#10 counter$count = 67068;
	#10 counter$count = 67069;
	#10 counter$count = 67070;
	#10 counter$count = 67071;
	#10 counter$count = 67072;
	#10 counter$count = 67073;
	#10 counter$count = 67074;
	#10 counter$count = 67075;
	#10 counter$count = 67076;
	#10 counter$count = 67077;
	#10 counter$count = 67078;
	#10 counter$count = 67079;
	#10 counter$count = 67080;
	#10 counter$count = 67081;
	#10 counter$count = 67082;
	#10 counter$count = 67083;
	#10 counter$count = 67084;
	#10 counter$count = 67085;
	#10 counter$count = 67086;
	#10 counter$count = 67087;
	#10 counter$count = 67088;
	#10 counter$count = 67089;
	#10 counter$count = 67090;
	#10 counter$count = 67091;
	#10 counter$count = 67092;
	#10 counter$count = 67093;
	#10 counter$count = 67094;
	#10 counter$count = 67095;
	#10 counter$count = 67096;
	#10 counter$count = 67097;
	#10 counter$count = 67098;
	#10 counter$count = 67099;
	#10 counter$count = 67100;
	#10 counter$count = 67101;
	#10 counter$count = 67102;
	#10 counter$count = 67103;
	#10 counter$count = 67104;
	#10 counter$count = 67105;
	#10 counter$count = 67106;
	#10 counter$count = 67107;
	#10 counter$count = 67108;
	#10 counter$count = 67109;
	#10 counter$count = 67110;
	#10 counter$count = 67111;
	#10 counter$count = 67112;
	#10 counter$count = 67113;
	#10 counter$count = 67114;
	#10 counter$count = 67115;
	#10 counter$count = 67116;
	#10 counter$count = 67117;
	#10 counter$count = 67118;
	#10 counter$count = 67119;
	#10 counter$count = 67120;
	#10 counter$count = 67121;
	#10 counter$count = 67122;
	#10 counter$count = 67123;
	#10 counter$count = 67124;
	#10 counter$count = 67125;
	#10 counter$count = 67126;
	#10 counter$count = 67127;
	#10 counter$count = 67128;
	#10 counter$count = 67129;
	#10 counter$count = 67130;
	#10 counter$count = 67131;
	#10 counter$count = 67132;
	#10 counter$count = 67133;
	#10 counter$count = 67134;
	#10 counter$count = 67135;
	#10 counter$count = 67136;
	#10 counter$count = 67137;
	#10 counter$count = 67138;
	#10 counter$count = 67139;
	#10 counter$count = 67140;
	#10 counter$count = 67141;
	#10 counter$count = 67142;
	#10 counter$count = 67143;
	#10 counter$count = 67144;
	#10 counter$count = 67145;
	#10 counter$count = 67146;
	#10 counter$count = 67147;
	#10 counter$count = 67148;
	#10 counter$count = 67149;
	#10 counter$count = 67150;
	#10 counter$count = 67151;
	#10 counter$count = 67152;
	#10 counter$count = 67153;
	#10 counter$count = 67154;
	#10 counter$count = 67155;
	#10 counter$count = 67156;
	#10 counter$count = 67157;
	#10 counter$count = 67158;
	#10 counter$count = 67159;
	#10 counter$count = 67160;
	#10 counter$count = 67161;
	#10 counter$count = 67162;
	#10 counter$count = 67163;
	#10 counter$count = 67164;
	#10 counter$count = 67165;
	#10 counter$count = 67166;
	#10 counter$count = 67167;
	#10 counter$count = 67168;
	#10 counter$count = 67169;
	#10 counter$count = 67170;
	#10 counter$count = 67171;
	#10 counter$count = 67172;
	#10 counter$count = 67173;
	#10 counter$count = 67174;
	#10 counter$count = 67175;
	#10 counter$count = 67176;
	#10 counter$count = 67177;
	#10 counter$count = 67178;
	#10 counter$count = 67179;
	#10 counter$count = 67180;
	#10 counter$count = 67181;
	#10 counter$count = 67182;
	#10 counter$count = 67183;
	#10 counter$count = 67184;
	#10 counter$count = 67185;
	#10 counter$count = 67186;
	#10 counter$count = 67187;
	#10 counter$count = 67188;
	#10 counter$count = 67189;
	#10 counter$count = 67190;
	#10 counter$count = 67191;
	#10 counter$count = 67192;
	#10 counter$count = 67193;
	#10 counter$count = 67194;
	#10 counter$count = 67195;
	#10 counter$count = 67196;
	#10 counter$count = 67197;
	#10 counter$count = 67198;
	#10 counter$count = 67199;
	#10 counter$count = 67200;
	#10 counter$count = 67201;
	#10 counter$count = 67202;
	#10 counter$count = 67203;
	#10 counter$count = 67204;
	#10 counter$count = 67205;
	#10 counter$count = 67206;
	#10 counter$count = 67207;
	#10 counter$count = 67208;
	#10 counter$count = 67209;
	#10 counter$count = 67210;
	#10 counter$count = 67211;
	#10 counter$count = 67212;
	#10 counter$count = 67213;
	#10 counter$count = 67214;
	#10 counter$count = 67215;
	#10 counter$count = 67216;
	#10 counter$count = 67217;
	#10 counter$count = 67218;
	#10 counter$count = 67219;
	#10 counter$count = 67220;
	#10 counter$count = 67221;
	#10 counter$count = 67222;
	#10 counter$count = 67223;
	#10 counter$count = 67224;
	#10 counter$count = 67225;
	#10 counter$count = 67226;
	#10 counter$count = 67227;
	#10 counter$count = 67228;
	#10 counter$count = 67229;
	#10 counter$count = 67230;
	#10 counter$count = 67231;
	#10 counter$count = 67232;
	#10 counter$count = 67233;
	#10 counter$count = 67234;
	#10 counter$count = 67235;
	#10 counter$count = 67236;
	#10 counter$count = 67237;
	#10 counter$count = 67238;
	#10 counter$count = 67239;
	#10 counter$count = 67240;
	#10 counter$count = 67241;
	#10 counter$count = 67242;
	#10 counter$count = 67243;
	#10 counter$count = 67244;
	#10 counter$count = 67245;
	#10 counter$count = 67246;
	#10 counter$count = 67247;
	#10 counter$count = 67248;
	#10 counter$count = 67249;
	#10 counter$count = 67250;
	#10 counter$count = 67251;
	#10 counter$count = 67252;
	#10 counter$count = 67253;
	#10 counter$count = 67254;
	#10 counter$count = 67255;
	#10 counter$count = 67256;
	#10 counter$count = 67257;
	#10 counter$count = 67258;
	#10 counter$count = 67259;
	#10 counter$count = 67260;
	#10 counter$count = 67261;
	#10 counter$count = 67262;
	#10 counter$count = 67263;
	#10 counter$count = 67264;
	#10 counter$count = 67265;
	#10 counter$count = 67266;
	#10 counter$count = 67267;
	#10 counter$count = 67268;
	#10 counter$count = 67269;
	#10 counter$count = 67270;
	#10 counter$count = 67271;
	#10 counter$count = 67272;
	#10 counter$count = 67273;
	#10 counter$count = 67274;
	#10 counter$count = 67275;
	#10 counter$count = 67276;
	#10 counter$count = 67277;
	#10 counter$count = 67278;
	#10 counter$count = 67279;
	#10 counter$count = 67280;
	#10 counter$count = 67281;
	#10 counter$count = 67282;
	#10 counter$count = 67283;
	#10 counter$count = 67284;
	#10 counter$count = 67285;
	#10 counter$count = 67286;
	#10 counter$count = 67287;
	#10 counter$count = 67288;
	#10 counter$count = 67289;
	#10 counter$count = 67290;
	#10 counter$count = 67291;
	#10 counter$count = 67292;
	#10 counter$count = 67293;
	#10 counter$count = 67294;
	#10 counter$count = 67295;
	#10 counter$count = 67296;
	#10 counter$count = 67297;
	#10 counter$count = 67298;
	#10 counter$count = 67299;
	#10 counter$count = 67300;
	#10 counter$count = 67301;
	#10 counter$count = 67302;
	#10 counter$count = 67303;
	#10 counter$count = 67304;
	#10 counter$count = 67305;
	#10 counter$count = 67306;
	#10 counter$count = 67307;
	#10 counter$count = 67308;
	#10 counter$count = 67309;
	#10 counter$count = 67310;
	#10 counter$count = 67311;
	#10 counter$count = 67312;
	#10 counter$count = 67313;
	#10 counter$count = 67314;
	#10 counter$count = 67315;
	#10 counter$count = 67316;
	#10 counter$count = 67317;
	#10 counter$count = 67318;
	#10 counter$count = 67319;
	#10 counter$count = 67320;
	#10 counter$count = 67321;
	#10 counter$count = 67322;
	#10 counter$count = 67323;
	#10 counter$count = 67324;
	#10 counter$count = 67325;
	#10 counter$count = 67326;
	#10 counter$count = 67327;
	#10 counter$count = 67328;
	#10 counter$count = 67329;
	#10 counter$count = 67330;
	#10 counter$count = 67331;
	#10 counter$count = 67332;
	#10 counter$count = 67333;
	#10 counter$count = 67334;
	#10 counter$count = 67335;
	#10 counter$count = 67336;
	#10 counter$count = 67337;
	#10 counter$count = 67338;
	#10 counter$count = 67339;
	#10 counter$count = 67340;
	#10 counter$count = 67341;
	#10 counter$count = 67342;
	#10 counter$count = 67343;
	#10 counter$count = 67344;
	#10 counter$count = 67345;
	#10 counter$count = 67346;
	#10 counter$count = 67347;
	#10 counter$count = 67348;
	#10 counter$count = 67349;
	#10 counter$count = 67350;
	#10 counter$count = 67351;
	#10 counter$count = 67352;
	#10 counter$count = 67353;
	#10 counter$count = 67354;
	#10 counter$count = 67355;
	#10 counter$count = 67356;
	#10 counter$count = 67357;
	#10 counter$count = 67358;
	#10 counter$count = 67359;
	#10 counter$count = 67360;
	#10 counter$count = 67361;
	#10 counter$count = 67362;
	#10 counter$count = 67363;
	#10 counter$count = 67364;
	#10 counter$count = 67365;
	#10 counter$count = 67366;
	#10 counter$count = 67367;
	#10 counter$count = 67368;
	#10 counter$count = 67369;
	#10 counter$count = 67370;
	#10 counter$count = 67371;
	#10 counter$count = 67372;
	#10 counter$count = 67373;
	#10 counter$count = 67374;
	#10 counter$count = 67375;
	#10 counter$count = 67376;
	#10 counter$count = 67377;
	#10 counter$count = 67378;
	#10 counter$count = 67379;
	#10 counter$count = 67380;
	#10 counter$count = 67381;
	#10 counter$count = 67382;
	#10 counter$count = 67383;
	#10 counter$count = 67384;
	#10 counter$count = 67385;
	#10 counter$count = 67386;
	#10 counter$count = 67387;
	#10 counter$count = 67388;
	#10 counter$count = 67389;
	#10 counter$count = 67390;
	#10 counter$count = 67391;
	#10 counter$count = 67392;
	#10 counter$count = 67393;
	#10 counter$count = 67394;
	#10 counter$count = 67395;
	#10 counter$count = 67396;
	#10 counter$count = 67397;
	#10 counter$count = 67398;
	#10 counter$count = 67399;
	#10 counter$count = 67400;
	#10 counter$count = 67401;
	#10 counter$count = 67402;
	#10 counter$count = 67403;
	#10 counter$count = 67404;
	#10 counter$count = 67405;
	#10 counter$count = 67406;
	#10 counter$count = 67407;
	#10 counter$count = 67408;
	#10 counter$count = 67409;
	#10 counter$count = 67410;
	#10 counter$count = 67411;
	#10 counter$count = 67412;
	#10 counter$count = 67413;
	#10 counter$count = 67414;
	#10 counter$count = 67415;
	#10 counter$count = 67416;
	#10 counter$count = 67417;
	#10 counter$count = 67418;
	#10 counter$count = 67419;
	#10 counter$count = 67420;
	#10 counter$count = 67421;
	#10 counter$count = 67422;
	#10 counter$count = 67423;
	#10 counter$count = 67424;
	#10 counter$count = 67425;
	#10 counter$count = 67426;
	#10 counter$count = 67427;
	#10 counter$count = 67428;
	#10 counter$count = 67429;
	#10 counter$count = 67430;
	#10 counter$count = 67431;
	#10 counter$count = 67432;
	#10 counter$count = 67433;
	#10 counter$count = 67434;
	#10 counter$count = 67435;
	#10 counter$count = 67436;
	#10 counter$count = 67437;
	#10 counter$count = 67438;
	#10 counter$count = 67439;
	#10 counter$count = 67440;
	#10 counter$count = 67441;
	#10 counter$count = 67442;
	#10 counter$count = 67443;
	#10 counter$count = 67444;
	#10 counter$count = 67445;
	#10 counter$count = 67446;
	#10 counter$count = 67447;
	#10 counter$count = 67448;
	#10 counter$count = 67449;
	#10 counter$count = 67450;
	#10 counter$count = 67451;
	#10 counter$count = 67452;
	#10 counter$count = 67453;
	#10 counter$count = 67454;
	#10 counter$count = 67455;
	#10 counter$count = 67456;
	#10 counter$count = 67457;
	#10 counter$count = 67458;
	#10 counter$count = 67459;
	#10 counter$count = 67460;
	#10 counter$count = 67461;
	#10 counter$count = 67462;
	#10 counter$count = 67463;
	#10 counter$count = 67464;
	#10 counter$count = 67465;
	#10 counter$count = 67466;
	#10 counter$count = 67467;
	#10 counter$count = 67468;
	#10 counter$count = 67469;
	#10 counter$count = 67470;
	#10 counter$count = 67471;
	#10 counter$count = 67472;
	#10 counter$count = 67473;
	#10 counter$count = 67474;
	#10 counter$count = 67475;
	#10 counter$count = 67476;
	#10 counter$count = 67477;
	#10 counter$count = 67478;
	#10 counter$count = 67479;
	#10 counter$count = 67480;
	#10 counter$count = 67481;
	#10 counter$count = 67482;
	#10 counter$count = 67483;
	#10 counter$count = 67484;
	#10 counter$count = 67485;
	#10 counter$count = 67486;
	#10 counter$count = 67487;
	#10 counter$count = 67488;
	#10 counter$count = 67489;
	#10 counter$count = 67490;
	#10 counter$count = 67491;
	#10 counter$count = 67492;
	#10 counter$count = 67493;
	#10 counter$count = 67494;
	#10 counter$count = 67495;
	#10 counter$count = 67496;
	#10 counter$count = 67497;
	#10 counter$count = 67498;
	#10 counter$count = 67499;
	#10 counter$count = 67500;
	#10 counter$count = 67501;
	#10 counter$count = 67502;
	#10 counter$count = 67503;
	#10 counter$count = 67504;
	#10 counter$count = 67505;
	#10 counter$count = 67506;
	#10 counter$count = 67507;
	#10 counter$count = 67508;
	#10 counter$count = 67509;
	#10 counter$count = 67510;
	#10 counter$count = 67511;
	#10 counter$count = 67512;
	#10 counter$count = 67513;
	#10 counter$count = 67514;
	#10 counter$count = 67515;
	#10 counter$count = 67516;
	#10 counter$count = 67517;
	#10 counter$count = 67518;
	#10 counter$count = 67519;
	#10 counter$count = 67520;
	#10 counter$count = 67521;
	#10 counter$count = 67522;
	#10 counter$count = 67523;
	#10 counter$count = 67524;
	#10 counter$count = 67525;
	#10 counter$count = 67526;
	#10 counter$count = 67527;
	#10 counter$count = 67528;
	#10 counter$count = 67529;
	#10 counter$count = 67530;
	#10 counter$count = 67531;
	#10 counter$count = 67532;
	#10 counter$count = 67533;
	#10 counter$count = 67534;
	#10 counter$count = 67535;
	#10 counter$count = 67536;
	#10 counter$count = 67537;
	#10 counter$count = 67538;
	#10 counter$count = 67539;
	#10 counter$count = 67540;
	#10 counter$count = 67541;
	#10 counter$count = 67542;
	#10 counter$count = 67543;
	#10 counter$count = 67544;
	#10 counter$count = 67545;
	#10 counter$count = 67546;
	#10 counter$count = 67547;
	#10 counter$count = 67548;
	#10 counter$count = 67549;
	#10 counter$count = 67550;
	#10 counter$count = 67551;
	#10 counter$count = 67552;
	#10 counter$count = 67553;
	#10 counter$count = 67554;
	#10 counter$count = 67555;
	#10 counter$count = 67556;
	#10 counter$count = 67557;
	#10 counter$count = 67558;
	#10 counter$count = 67559;
	#10 counter$count = 67560;
	#10 counter$count = 67561;
	#10 counter$count = 67562;
	#10 counter$count = 67563;
	#10 counter$count = 67564;
	#10 counter$count = 67565;
	#10 counter$count = 67566;
	#10 counter$count = 67567;
	#10 counter$count = 67568;
	#10 counter$count = 67569;
	#10 counter$count = 67570;
	#10 counter$count = 67571;
	#10 counter$count = 67572;
	#10 counter$count = 67573;
	#10 counter$count = 67574;
	#10 counter$count = 67575;
	#10 counter$count = 67576;
	#10 counter$count = 67577;
	#10 counter$count = 67578;
	#10 counter$count = 67579;
	#10 counter$count = 67580;
	#10 counter$count = 67581;
	#10 counter$count = 67582;
	#10 counter$count = 67583;
	#10 counter$count = 67584;
	#10 counter$count = 67585;
	#10 counter$count = 67586;
	#10 counter$count = 67587;
	#10 counter$count = 67588;
	#10 counter$count = 67589;
	#10 counter$count = 67590;
	#10 counter$count = 67591;
	#10 counter$count = 67592;
	#10 counter$count = 67593;
	#10 counter$count = 67594;
	#10 counter$count = 67595;
	#10 counter$count = 67596;
	#10 counter$count = 67597;
	#10 counter$count = 67598;
	#10 counter$count = 67599;
	#10 counter$count = 67600;
	#10 counter$count = 67601;
	#10 counter$count = 67602;
	#10 counter$count = 67603;
	#10 counter$count = 67604;
	#10 counter$count = 67605;
	#10 counter$count = 67606;
	#10 counter$count = 67607;
	#10 counter$count = 67608;
	#10 counter$count = 67609;
	#10 counter$count = 67610;
	#10 counter$count = 67611;
	#10 counter$count = 67612;
	#10 counter$count = 67613;
	#10 counter$count = 67614;
	#10 counter$count = 67615;
	#10 counter$count = 67616;
	#10 counter$count = 67617;
	#10 counter$count = 67618;
	#10 counter$count = 67619;
	#10 counter$count = 67620;
	#10 counter$count = 67621;
	#10 counter$count = 67622;
	#10 counter$count = 67623;
	#10 counter$count = 67624;
	#10 counter$count = 67625;
	#10 counter$count = 67626;
	#10 counter$count = 67627;
	#10 counter$count = 67628;
	#10 counter$count = 67629;
	#10 counter$count = 67630;
	#10 counter$count = 67631;
	#10 counter$count = 67632;
	#10 counter$count = 67633;
	#10 counter$count = 67634;
	#10 counter$count = 67635;
	#10 counter$count = 67636;
	#10 counter$count = 67637;
	#10 counter$count = 67638;
	#10 counter$count = 67639;
	#10 counter$count = 67640;
	#10 counter$count = 67641;
	#10 counter$count = 67642;
	#10 counter$count = 67643;
	#10 counter$count = 67644;
	#10 counter$count = 67645;
	#10 counter$count = 67646;
	#10 counter$count = 67647;
	#10 counter$count = 67648;
	#10 counter$count = 67649;
	#10 counter$count = 67650;
	#10 counter$count = 67651;
	#10 counter$count = 67652;
	#10 counter$count = 67653;
	#10 counter$count = 67654;
	#10 counter$count = 67655;
	#10 counter$count = 67656;
	#10 counter$count = 67657;
	#10 counter$count = 67658;
	#10 counter$count = 67659;
	#10 counter$count = 67660;
	#10 counter$count = 67661;
	#10 counter$count = 67662;
	#10 counter$count = 67663;
	#10 counter$count = 67664;
	#10 counter$count = 67665;
	#10 counter$count = 67666;
	#10 counter$count = 67667;
	#10 counter$count = 67668;
	#10 counter$count = 67669;
	#10 counter$count = 67670;
	#10 counter$count = 67671;
	#10 counter$count = 67672;
	#10 counter$count = 67673;
	#10 counter$count = 67674;
	#10 counter$count = 67675;
	#10 counter$count = 67676;
	#10 counter$count = 67677;
	#10 counter$count = 67678;
	#10 counter$count = 67679;
	#10 counter$count = 67680;
	#10 counter$count = 67681;
	#10 counter$count = 67682;
	#10 counter$count = 67683;
	#10 counter$count = 67684;
	#10 counter$count = 67685;
	#10 counter$count = 67686;
	#10 counter$count = 67687;
	#10 counter$count = 67688;
	#10 counter$count = 67689;
	#10 counter$count = 67690;
	#10 counter$count = 67691;
	#10 counter$count = 67692;
	#10 counter$count = 67693;
	#10 counter$count = 67694;
	#10 counter$count = 67695;
	#10 counter$count = 67696;
	#10 counter$count = 67697;
	#10 counter$count = 67698;
	#10 counter$count = 67699;
	#10 counter$count = 67700;
	#10 counter$count = 67701;
	#10 counter$count = 67702;
	#10 counter$count = 67703;
	#10 counter$count = 67704;
	#10 counter$count = 67705;
	#10 counter$count = 67706;
	#10 counter$count = 67707;
	#10 counter$count = 67708;
	#10 counter$count = 67709;
	#10 counter$count = 67710;
	#10 counter$count = 67711;
	#10 counter$count = 67712;
	#10 counter$count = 67713;
	#10 counter$count = 67714;
	#10 counter$count = 67715;
	#10 counter$count = 67716;
	#10 counter$count = 67717;
	#10 counter$count = 67718;
	#10 counter$count = 67719;
	#10 counter$count = 67720;
	#10 counter$count = 67721;
	#10 counter$count = 67722;
	#10 counter$count = 67723;
	#10 counter$count = 67724;
	#10 counter$count = 67725;
	#10 counter$count = 67726;
	#10 counter$count = 67727;
	#10 counter$count = 67728;
	#10 counter$count = 67729;
	#10 counter$count = 67730;
	#10 counter$count = 67731;
	#10 counter$count = 67732;
	#10 counter$count = 67733;
	#10 counter$count = 67734;
	#10 counter$count = 67735;
	#10 counter$count = 67736;
	#10 counter$count = 67737;
	#10 counter$count = 67738;
	#10 counter$count = 67739;
	#10 counter$count = 67740;
	#10 counter$count = 67741;
	#10 counter$count = 67742;
	#10 counter$count = 67743;
	#10 counter$count = 67744;
	#10 counter$count = 67745;
	#10 counter$count = 67746;
	#10 counter$count = 67747;
	#10 counter$count = 67748;
	#10 counter$count = 67749;
	#10 counter$count = 67750;
	#10 counter$count = 67751;
	#10 counter$count = 67752;
	#10 counter$count = 67753;
	#10 counter$count = 67754;
	#10 counter$count = 67755;
	#10 counter$count = 67756;
	#10 counter$count = 67757;
	#10 counter$count = 67758;
	#10 counter$count = 67759;
	#10 counter$count = 67760;
	#10 counter$count = 67761;
	#10 counter$count = 67762;
	#10 counter$count = 67763;
	#10 counter$count = 67764;
	#10 counter$count = 67765;
	#10 counter$count = 67766;
	#10 counter$count = 67767;
	#10 counter$count = 67768;
	#10 counter$count = 67769;
	#10 counter$count = 67770;
	#10 counter$count = 67771;
	#10 counter$count = 67772;
	#10 counter$count = 67773;
	#10 counter$count = 67774;
	#10 counter$count = 67775;
	#10 counter$count = 67776;
	#10 counter$count = 67777;
	#10 counter$count = 67778;
	#10 counter$count = 67779;
	#10 counter$count = 67780;
	#10 counter$count = 67781;
	#10 counter$count = 67782;
	#10 counter$count = 67783;
	#10 counter$count = 67784;
	#10 counter$count = 67785;
	#10 counter$count = 67786;
	#10 counter$count = 67787;
	#10 counter$count = 67788;
	#10 counter$count = 67789;
	#10 counter$count = 67790;
	#10 counter$count = 67791;
	#10 counter$count = 67792;
	#10 counter$count = 67793;
	#10 counter$count = 67794;
	#10 counter$count = 67795;
	#10 counter$count = 67796;
	#10 counter$count = 67797;
	#10 counter$count = 67798;
	#10 counter$count = 67799;
	#10 counter$count = 67800;
	#10 counter$count = 67801;
	#10 counter$count = 67802;
	#10 counter$count = 67803;
	#10 counter$count = 67804;
	#10 counter$count = 67805;
	#10 counter$count = 67806;
	#10 counter$count = 67807;
	#10 counter$count = 67808;
	#10 counter$count = 67809;
	#10 counter$count = 67810;
	#10 counter$count = 67811;
	#10 counter$count = 67812;
	#10 counter$count = 67813;
	#10 counter$count = 67814;
	#10 counter$count = 67815;
	#10 counter$count = 67816;
	#10 counter$count = 67817;
	#10 counter$count = 67818;
	#10 counter$count = 67819;
	#10 counter$count = 67820;
	#10 counter$count = 67821;
	#10 counter$count = 67822;
	#10 counter$count = 67823;
	#10 counter$count = 67824;
	#10 counter$count = 67825;
	#10 counter$count = 67826;
	#10 counter$count = 67827;
	#10 counter$count = 67828;
	#10 counter$count = 67829;
	#10 counter$count = 67830;
	#10 counter$count = 67831;
	#10 counter$count = 67832;
	#10 counter$count = 67833;
	#10 counter$count = 67834;
	#10 counter$count = 67835;
	#10 counter$count = 67836;
	#10 counter$count = 67837;
	#10 counter$count = 67838;
	#10 counter$count = 67839;
	#10 counter$count = 67840;
	#10 counter$count = 67841;
	#10 counter$count = 67842;
	#10 counter$count = 67843;
	#10 counter$count = 67844;
	#10 counter$count = 67845;
	#10 counter$count = 67846;
	#10 counter$count = 67847;
	#10 counter$count = 67848;
	#10 counter$count = 67849;
	#10 counter$count = 67850;
	#10 counter$count = 67851;
	#10 counter$count = 67852;
	#10 counter$count = 67853;
	#10 counter$count = 67854;
	#10 counter$count = 67855;
	#10 counter$count = 67856;
	#10 counter$count = 67857;
	#10 counter$count = 67858;
	#10 counter$count = 67859;
	#10 counter$count = 67860;
	#10 counter$count = 67861;
	#10 counter$count = 67862;
	#10 counter$count = 67863;
	#10 counter$count = 67864;
	#10 counter$count = 67865;
	#10 counter$count = 67866;
	#10 counter$count = 67867;
	#10 counter$count = 67868;
	#10 counter$count = 67869;
	#10 counter$count = 67870;
	#10 counter$count = 67871;
	#10 counter$count = 67872;
	#10 counter$count = 67873;
	#10 counter$count = 67874;
	#10 counter$count = 67875;
	#10 counter$count = 67876;
	#10 counter$count = 67877;
	#10 counter$count = 67878;
	#10 counter$count = 67879;
	#10 counter$count = 67880;
	#10 counter$count = 67881;
	#10 counter$count = 67882;
	#10 counter$count = 67883;
	#10 counter$count = 67884;
	#10 counter$count = 67885;
	#10 counter$count = 67886;
	#10 counter$count = 67887;
	#10 counter$count = 67888;
	#10 counter$count = 67889;
	#10 counter$count = 67890;
	#10 counter$count = 67891;
	#10 counter$count = 67892;
	#10 counter$count = 67893;
	#10 counter$count = 67894;
	#10 counter$count = 67895;
	#10 counter$count = 67896;
	#10 counter$count = 67897;
	#10 counter$count = 67898;
	#10 counter$count = 67899;
	#10 counter$count = 67900;
	#10 counter$count = 67901;
	#10 counter$count = 67902;
	#10 counter$count = 67903;
	#10 counter$count = 67904;
	#10 counter$count = 67905;
	#10 counter$count = 67906;
	#10 counter$count = 67907;
	#10 counter$count = 67908;
	#10 counter$count = 67909;
	#10 counter$count = 67910;
	#10 counter$count = 67911;
	#10 counter$count = 67912;
	#10 counter$count = 67913;
	#10 counter$count = 67914;
	#10 counter$count = 67915;
	#10 counter$count = 67916;
	#10 counter$count = 67917;
	#10 counter$count = 67918;
	#10 counter$count = 67919;
	#10 counter$count = 67920;
	#10 counter$count = 67921;
	#10 counter$count = 67922;
	#10 counter$count = 67923;
	#10 counter$count = 67924;
	#10 counter$count = 67925;
	#10 counter$count = 67926;
	#10 counter$count = 67927;
	#10 counter$count = 67928;
	#10 counter$count = 67929;
	#10 counter$count = 67930;
	#10 counter$count = 67931;
	#10 counter$count = 67932;
	#10 counter$count = 67933;
	#10 counter$count = 67934;
	#10 counter$count = 67935;
	#10 counter$count = 67936;
	#10 counter$count = 67937;
	#10 counter$count = 67938;
	#10 counter$count = 67939;
	#10 counter$count = 67940;
	#10 counter$count = 67941;
	#10 counter$count = 67942;
	#10 counter$count = 67943;
	#10 counter$count = 67944;
	#10 counter$count = 67945;
	#10 counter$count = 67946;
	#10 counter$count = 67947;
	#10 counter$count = 67948;
	#10 counter$count = 67949;
	#10 counter$count = 67950;
	#10 counter$count = 67951;
	#10 counter$count = 67952;
	#10 counter$count = 67953;
	#10 counter$count = 67954;
	#10 counter$count = 67955;
	#10 counter$count = 67956;
	#10 counter$count = 67957;
	#10 counter$count = 67958;
	#10 counter$count = 67959;
	#10 counter$count = 67960;
	#10 counter$count = 67961;
	#10 counter$count = 67962;
	#10 counter$count = 67963;
	#10 counter$count = 67964;
	#10 counter$count = 67965;
	#10 counter$count = 67966;
	#10 counter$count = 67967;
	#10 counter$count = 67968;
	#10 counter$count = 67969;
	#10 counter$count = 67970;
	#10 counter$count = 67971;
	#10 counter$count = 67972;
	#10 counter$count = 67973;
	#10 counter$count = 67974;
	#10 counter$count = 67975;
	#10 counter$count = 67976;
	#10 counter$count = 67977;
	#10 counter$count = 67978;
	#10 counter$count = 67979;
	#10 counter$count = 67980;
	#10 counter$count = 67981;
	#10 counter$count = 67982;
	#10 counter$count = 67983;
	#10 counter$count = 67984;
	#10 counter$count = 67985;
	#10 counter$count = 67986;
	#10 counter$count = 67987;
	#10 counter$count = 67988;
	#10 counter$count = 67989;
	#10 counter$count = 67990;
	#10 counter$count = 67991;
	#10 counter$count = 67992;
	#10 counter$count = 67993;
	#10 counter$count = 67994;
	#10 counter$count = 67995;
	#10 counter$count = 67996;
	#10 counter$count = 67997;
	#10 counter$count = 67998;
	#10 counter$count = 67999;
	#10 counter$count = 68000;
	#10 counter$count = 68001;
	#10 counter$count = 68002;
	#10 counter$count = 68003;
	#10 counter$count = 68004;
	#10 counter$count = 68005;
	#10 counter$count = 68006;
	#10 counter$count = 68007;
	#10 counter$count = 68008;
	#10 counter$count = 68009;
	#10 counter$count = 68010;
	#10 counter$count = 68011;
	#10 counter$count = 68012;
	#10 counter$count = 68013;
	#10 counter$count = 68014;
	#10 counter$count = 68015;
	#10 counter$count = 68016;
	#10 counter$count = 68017;
	#10 counter$count = 68018;
	#10 counter$count = 68019;
	#10 counter$count = 68020;
	#10 counter$count = 68021;
	#10 counter$count = 68022;
	#10 counter$count = 68023;
	#10 counter$count = 68024;
	#10 counter$count = 68025;
	#10 counter$count = 68026;
	#10 counter$count = 68027;
	#10 counter$count = 68028;
	#10 counter$count = 68029;
	#10 counter$count = 68030;
	#10 counter$count = 68031;
	#10 counter$count = 68032;
	#10 counter$count = 68033;
	#10 counter$count = 68034;
	#10 counter$count = 68035;
	#10 counter$count = 68036;
	#10 counter$count = 68037;
	#10 counter$count = 68038;
	#10 counter$count = 68039;
	#10 counter$count = 68040;
	#10 counter$count = 68041;
	#10 counter$count = 68042;
	#10 counter$count = 68043;
	#10 counter$count = 68044;
	#10 counter$count = 68045;
	#10 counter$count = 68046;
	#10 counter$count = 68047;
	#10 counter$count = 68048;
	#10 counter$count = 68049;
	#10 counter$count = 68050;
	#10 counter$count = 68051;
	#10 counter$count = 68052;
	#10 counter$count = 68053;
	#10 counter$count = 68054;
	#10 counter$count = 68055;
	#10 counter$count = 68056;
	#10 counter$count = 68057;
	#10 counter$count = 68058;
	#10 counter$count = 68059;
	#10 counter$count = 68060;
	#10 counter$count = 68061;
	#10 counter$count = 68062;
	#10 counter$count = 68063;
	#10 counter$count = 68064;
	#10 counter$count = 68065;
	#10 counter$count = 68066;
	#10 counter$count = 68067;
	#10 counter$count = 68068;
	#10 counter$count = 68069;
	#10 counter$count = 68070;
	#10 counter$count = 68071;
	#10 counter$count = 68072;
	#10 counter$count = 68073;
	#10 counter$count = 68074;
	#10 counter$count = 68075;
	#10 counter$count = 68076;
	#10 counter$count = 68077;
	#10 counter$count = 68078;
	#10 counter$count = 68079;
	#10 counter$count = 68080;
	#10 counter$count = 68081;
	#10 counter$count = 68082;
	#10 counter$count = 68083;
	#10 counter$count = 68084;
	#10 counter$count = 68085;
	#10 counter$count = 68086;
	#10 counter$count = 68087;
	#10 counter$count = 68088;
	#10 counter$count = 68089;
	#10 counter$count = 68090;
	#10 counter$count = 68091;
	#10 counter$count = 68092;
	#10 counter$count = 68093;
	#10 counter$count = 68094;
	#10 counter$count = 68095;
	#10 counter$count = 68096;
	#10 counter$count = 68097;
	#10 counter$count = 68098;
	#10 counter$count = 68099;
	#10 counter$count = 68100;
	#10 counter$count = 68101;
	#10 counter$count = 68102;
	#10 counter$count = 68103;
	#10 counter$count = 68104;
	#10 counter$count = 68105;
	#10 counter$count = 68106;
	#10 counter$count = 68107;
	#10 counter$count = 68108;
	#10 counter$count = 68109;
	#10 counter$count = 68110;
	#10 counter$count = 68111;
	#10 counter$count = 68112;
	#10 counter$count = 68113;
	#10 counter$count = 68114;
	#10 counter$count = 68115;
	#10 counter$count = 68116;
	#10 counter$count = 68117;
	#10 counter$count = 68118;
	#10 counter$count = 68119;
	#10 counter$count = 68120;
	#10 counter$count = 68121;
	#10 counter$count = 68122;
	#10 counter$count = 68123;
	#10 counter$count = 68124;
	#10 counter$count = 68125;
	#10 counter$count = 68126;
	#10 counter$count = 68127;
	#10 counter$count = 68128;
	#10 counter$count = 68129;
	#10 counter$count = 68130;
	#10 counter$count = 68131;
	#10 counter$count = 68132;
	#10 counter$count = 68133;
	#10 counter$count = 68134;
	#10 counter$count = 68135;
	#10 counter$count = 68136;
	#10 counter$count = 68137;
	#10 counter$count = 68138;
	#10 counter$count = 68139;
	#10 counter$count = 68140;
	#10 counter$count = 68141;
	#10 counter$count = 68142;
	#10 counter$count = 68143;
	#10 counter$count = 68144;
	#10 counter$count = 68145;
	#10 counter$count = 68146;
	#10 counter$count = 68147;
	#10 counter$count = 68148;
	#10 counter$count = 68149;
	#10 counter$count = 68150;
	#10 counter$count = 68151;
	#10 counter$count = 68152;
	#10 counter$count = 68153;
	#10 counter$count = 68154;
	#10 counter$count = 68155;
	#10 counter$count = 68156;
	#10 counter$count = 68157;
	#10 counter$count = 68158;
	#10 counter$count = 68159;
	#10 counter$count = 68160;
	#10 counter$count = 68161;
	#10 counter$count = 68162;
	#10 counter$count = 68163;
	#10 counter$count = 68164;
	#10 counter$count = 68165;
	#10 counter$count = 68166;
	#10 counter$count = 68167;
	#10 counter$count = 68168;
	#10 counter$count = 68169;
	#10 counter$count = 68170;
	#10 counter$count = 68171;
	#10 counter$count = 68172;
	#10 counter$count = 68173;
	#10 counter$count = 68174;
	#10 counter$count = 68175;
	#10 counter$count = 68176;
	#10 counter$count = 68177;
	#10 counter$count = 68178;
	#10 counter$count = 68179;
	#10 counter$count = 68180;
	#10 counter$count = 68181;
	#10 counter$count = 68182;
	#10 counter$count = 68183;
	#10 counter$count = 68184;
	#10 counter$count = 68185;
	#10 counter$count = 68186;
	#10 counter$count = 68187;
	#10 counter$count = 68188;
	#10 counter$count = 68189;
	#10 counter$count = 68190;
	#10 counter$count = 68191;
	#10 counter$count = 68192;
	#10 counter$count = 68193;
	#10 counter$count = 68194;
	#10 counter$count = 68195;
	#10 counter$count = 68196;
	#10 counter$count = 68197;
	#10 counter$count = 68198;
	#10 counter$count = 68199;
	#10 counter$count = 68200;
	#10 counter$count = 68201;
	#10 counter$count = 68202;
	#10 counter$count = 68203;
	#10 counter$count = 68204;
	#10 counter$count = 68205;
	#10 counter$count = 68206;
	#10 counter$count = 68207;
	#10 counter$count = 68208;
	#10 counter$count = 68209;
	#10 counter$count = 68210;
	#10 counter$count = 68211;
	#10 counter$count = 68212;
	#10 counter$count = 68213;
	#10 counter$count = 68214;
	#10 counter$count = 68215;
	#10 counter$count = 68216;
	#10 counter$count = 68217;
	#10 counter$count = 68218;
	#10 counter$count = 68219;
	#10 counter$count = 68220;
	#10 counter$count = 68221;
	#10 counter$count = 68222;
	#10 counter$count = 68223;
	#10 counter$count = 68224;
	#10 counter$count = 68225;
	#10 counter$count = 68226;
	#10 counter$count = 68227;
	#10 counter$count = 68228;
	#10 counter$count = 68229;
	#10 counter$count = 68230;
	#10 counter$count = 68231;
	#10 counter$count = 68232;
	#10 counter$count = 68233;
	#10 counter$count = 68234;
	#10 counter$count = 68235;
	#10 counter$count = 68236;
	#10 counter$count = 68237;
	#10 counter$count = 68238;
	#10 counter$count = 68239;
	#10 counter$count = 68240;
	#10 counter$count = 68241;
	#10 counter$count = 68242;
	#10 counter$count = 68243;
	#10 counter$count = 68244;
	#10 counter$count = 68245;
	#10 counter$count = 68246;
	#10 counter$count = 68247;
	#10 counter$count = 68248;
	#10 counter$count = 68249;
	#10 counter$count = 68250;
	#10 counter$count = 68251;
	#10 counter$count = 68252;
	#10 counter$count = 68253;
	#10 counter$count = 68254;
	#10 counter$count = 68255;
	#10 counter$count = 68256;
	#10 counter$count = 68257;
	#10 counter$count = 68258;
	#10 counter$count = 68259;
	#10 counter$count = 68260;
	#10 counter$count = 68261;
	#10 counter$count = 68262;
	#10 counter$count = 68263;
	#10 counter$count = 68264;
	#10 counter$count = 68265;
	#10 counter$count = 68266;
	#10 counter$count = 68267;
	#10 counter$count = 68268;
	#10 counter$count = 68269;
	#10 counter$count = 68270;
	#10 counter$count = 68271;
	#10 counter$count = 68272;
	#10 counter$count = 68273;
	#10 counter$count = 68274;
	#10 counter$count = 68275;
	#10 counter$count = 68276;
	#10 counter$count = 68277;
	#10 counter$count = 68278;
	#10 counter$count = 68279;
	#10 counter$count = 68280;
	#10 counter$count = 68281;
	#10 counter$count = 68282;
	#10 counter$count = 68283;
	#10 counter$count = 68284;
	#10 counter$count = 68285;
	#10 counter$count = 68286;
	#10 counter$count = 68287;
	#10 counter$count = 68288;
	#10 counter$count = 68289;
	#10 counter$count = 68290;
	#10 counter$count = 68291;
	#10 counter$count = 68292;
	#10 counter$count = 68293;
	#10 counter$count = 68294;
	#10 counter$count = 68295;
	#10 counter$count = 68296;
	#10 counter$count = 68297;
	#10 counter$count = 68298;
	#10 counter$count = 68299;
	#10 counter$count = 68300;
	#10 counter$count = 68301;
	#10 counter$count = 68302;
	#10 counter$count = 68303;
	#10 counter$count = 68304;
	#10 counter$count = 68305;
	#10 counter$count = 68306;
	#10 counter$count = 68307;
	#10 counter$count = 68308;
	#10 counter$count = 68309;
	#10 counter$count = 68310;
	#10 counter$count = 68311;
	#10 counter$count = 68312;
	#10 counter$count = 68313;
	#10 counter$count = 68314;
	#10 counter$count = 68315;
	#10 counter$count = 68316;
	#10 counter$count = 68317;
	#10 counter$count = 68318;
	#10 counter$count = 68319;
	#10 counter$count = 68320;
	#10 counter$count = 68321;
	#10 counter$count = 68322;
	#10 counter$count = 68323;
	#10 counter$count = 68324;
	#10 counter$count = 68325;
	#10 counter$count = 68326;
	#10 counter$count = 68327;
	#10 counter$count = 68328;
	#10 counter$count = 68329;
	#10 counter$count = 68330;
	#10 counter$count = 68331;
	#10 counter$count = 68332;
	#10 counter$count = 68333;
	#10 counter$count = 68334;
	#10 counter$count = 68335;
	#10 counter$count = 68336;
	#10 counter$count = 68337;
	#10 counter$count = 68338;
	#10 counter$count = 68339;
	#10 counter$count = 68340;
	#10 counter$count = 68341;
	#10 counter$count = 68342;
	#10 counter$count = 68343;
	#10 counter$count = 68344;
	#10 counter$count = 68345;
	#10 counter$count = 68346;
	#10 counter$count = 68347;
	#10 counter$count = 68348;
	#10 counter$count = 68349;
	#10 counter$count = 68350;
	#10 counter$count = 68351;
	#10 counter$count = 68352;
	#10 counter$count = 68353;
	#10 counter$count = 68354;
	#10 counter$count = 68355;
	#10 counter$count = 68356;
	#10 counter$count = 68357;
	#10 counter$count = 68358;
	#10 counter$count = 68359;
	#10 counter$count = 68360;
	#10 counter$count = 68361;
	#10 counter$count = 68362;
	#10 counter$count = 68363;
	#10 counter$count = 68364;
	#10 counter$count = 68365;
	#10 counter$count = 68366;
	#10 counter$count = 68367;
	#10 counter$count = 68368;
	#10 counter$count = 68369;
	#10 counter$count = 68370;
	#10 counter$count = 68371;
	#10 counter$count = 68372;
	#10 counter$count = 68373;
	#10 counter$count = 68374;
	#10 counter$count = 68375;
	#10 counter$count = 68376;
	#10 counter$count = 68377;
	#10 counter$count = 68378;
	#10 counter$count = 68379;
	#10 counter$count = 68380;
	#10 counter$count = 68381;
	#10 counter$count = 68382;
	#10 counter$count = 68383;
	#10 counter$count = 68384;
	#10 counter$count = 68385;
	#10 counter$count = 68386;
	#10 counter$count = 68387;
	#10 counter$count = 68388;
	#10 counter$count = 68389;
	#10 counter$count = 68390;
	#10 counter$count = 68391;
	#10 counter$count = 68392;
	#10 counter$count = 68393;
	#10 counter$count = 68394;
	#10 counter$count = 68395;
	#10 counter$count = 68396;
	#10 counter$count = 68397;
	#10 counter$count = 68398;
	#10 counter$count = 68399;
	#10 counter$count = 68400;
	#10 counter$count = 68401;
	#10 counter$count = 68402;
	#10 counter$count = 68403;
	#10 counter$count = 68404;
	#10 counter$count = 68405;
	#10 counter$count = 68406;
	#10 counter$count = 68407;
	#10 counter$count = 68408;
	#10 counter$count = 68409;
	#10 counter$count = 68410;
	#10 counter$count = 68411;
	#10 counter$count = 68412;
	#10 counter$count = 68413;
	#10 counter$count = 68414;
	#10 counter$count = 68415;
	#10 counter$count = 68416;
	#10 counter$count = 68417;
	#10 counter$count = 68418;
	#10 counter$count = 68419;
	#10 counter$count = 68420;
	#10 counter$count = 68421;
	#10 counter$count = 68422;
	#10 counter$count = 68423;
	#10 counter$count = 68424;
	#10 counter$count = 68425;
	#10 counter$count = 68426;
	#10 counter$count = 68427;
	#10 counter$count = 68428;
	#10 counter$count = 68429;
	#10 counter$count = 68430;
	#10 counter$count = 68431;
	#10 counter$count = 68432;
	#10 counter$count = 68433;
	#10 counter$count = 68434;
	#10 counter$count = 68435;
	#10 counter$count = 68436;
	#10 counter$count = 68437;
	#10 counter$count = 68438;
	#10 counter$count = 68439;
	#10 counter$count = 68440;
	#10 counter$count = 68441;
	#10 counter$count = 68442;
	#10 counter$count = 68443;
	#10 counter$count = 68444;
	#10 counter$count = 68445;
	#10 counter$count = 68446;
	#10 counter$count = 68447;
	#10 counter$count = 68448;
	#10 counter$count = 68449;
	#10 counter$count = 68450;
	#10 counter$count = 68451;
	#10 counter$count = 68452;
	#10 counter$count = 68453;
	#10 counter$count = 68454;
	#10 counter$count = 68455;
	#10 counter$count = 68456;
	#10 counter$count = 68457;
	#10 counter$count = 68458;
	#10 counter$count = 68459;
	#10 counter$count = 68460;
	#10 counter$count = 68461;
	#10 counter$count = 68462;
	#10 counter$count = 68463;
	#10 counter$count = 68464;
	#10 counter$count = 68465;
	#10 counter$count = 68466;
	#10 counter$count = 68467;
	#10 counter$count = 68468;
	#10 counter$count = 68469;
	#10 counter$count = 68470;
	#10 counter$count = 68471;
	#10 counter$count = 68472;
	#10 counter$count = 68473;
	#10 counter$count = 68474;
	#10 counter$count = 68475;
	#10 counter$count = 68476;
	#10 counter$count = 68477;
	#10 counter$count = 68478;
	#10 counter$count = 68479;
	#10 counter$count = 68480;
	#10 counter$count = 68481;
	#10 counter$count = 68482;
	#10 counter$count = 68483;
	#10 counter$count = 68484;
	#10 counter$count = 68485;
	#10 counter$count = 68486;
	#10 counter$count = 68487;
	#10 counter$count = 68488;
	#10 counter$count = 68489;
	#10 counter$count = 68490;
	#10 counter$count = 68491;
	#10 counter$count = 68492;
	#10 counter$count = 68493;
	#10 counter$count = 68494;
	#10 counter$count = 68495;
	#10 counter$count = 68496;
	#10 counter$count = 68497;
	#10 counter$count = 68498;
	#10 counter$count = 68499;
	#10 counter$count = 68500;
	#10 counter$count = 68501;
	#10 counter$count = 68502;
	#10 counter$count = 68503;
	#10 counter$count = 68504;
	#10 counter$count = 68505;
	#10 counter$count = 68506;
	#10 counter$count = 68507;
	#10 counter$count = 68508;
	#10 counter$count = 68509;
	#10 counter$count = 68510;
	#10 counter$count = 68511;
	#10 counter$count = 68512;
	#10 counter$count = 68513;
	#10 counter$count = 68514;
	#10 counter$count = 68515;
	#10 counter$count = 68516;
	#10 counter$count = 68517;
	#10 counter$count = 68518;
	#10 counter$count = 68519;
	#10 counter$count = 68520;
	#10 counter$count = 68521;
	#10 counter$count = 68522;
	#10 counter$count = 68523;
	#10 counter$count = 68524;
	#10 counter$count = 68525;
	#10 counter$count = 68526;
	#10 counter$count = 68527;
	#10 counter$count = 68528;
	#10 counter$count = 68529;
	#10 counter$count = 68530;
	#10 counter$count = 68531;
	#10 counter$count = 68532;
	#10 counter$count = 68533;
	#10 counter$count = 68534;
	#10 counter$count = 68535;
	#10 counter$count = 68536;
	#10 counter$count = 68537;
	#10 counter$count = 68538;
	#10 counter$count = 68539;
	#10 counter$count = 68540;
	#10 counter$count = 68541;
	#10 counter$count = 68542;
	#10 counter$count = 68543;
	#10 counter$count = 68544;
	#10 counter$count = 68545;
	#10 counter$count = 68546;
	#10 counter$count = 68547;
	#10 counter$count = 68548;
	#10 counter$count = 68549;
	#10 counter$count = 68550;
	#10 counter$count = 68551;
	#10 counter$count = 68552;
	#10 counter$count = 68553;
	#10 counter$count = 68554;
	#10 counter$count = 68555;
	#10 counter$count = 68556;
	#10 counter$count = 68557;
	#10 counter$count = 68558;
	#10 counter$count = 68559;
	#10 counter$count = 68560;
	#10 counter$count = 68561;
	#10 counter$count = 68562;
	#10 counter$count = 68563;
	#10 counter$count = 68564;
	#10 counter$count = 68565;
	#10 counter$count = 68566;
	#10 counter$count = 68567;
	#10 counter$count = 68568;
	#10 counter$count = 68569;
	#10 counter$count = 68570;
	#10 counter$count = 68571;
	#10 counter$count = 68572;
	#10 counter$count = 68573;
	#10 counter$count = 68574;
	#10 counter$count = 68575;
	#10 counter$count = 68576;
	#10 counter$count = 68577;
	#10 counter$count = 68578;
	#10 counter$count = 68579;
	#10 counter$count = 68580;
	#10 counter$count = 68581;
	#10 counter$count = 68582;
	#10 counter$count = 68583;
	#10 counter$count = 68584;
	#10 counter$count = 68585;
	#10 counter$count = 68586;
	#10 counter$count = 68587;
	#10 counter$count = 68588;
	#10 counter$count = 68589;
	#10 counter$count = 68590;
	#10 counter$count = 68591;
	#10 counter$count = 68592;
	#10 counter$count = 68593;
	#10 counter$count = 68594;
	#10 counter$count = 68595;
	#10 counter$count = 68596;
	#10 counter$count = 68597;
	#10 counter$count = 68598;
	#10 counter$count = 68599;
	#10 counter$count = 68600;
	#10 counter$count = 68601;
	#10 counter$count = 68602;
	#10 counter$count = 68603;
	#10 counter$count = 68604;
	#10 counter$count = 68605;
	#10 counter$count = 68606;
	#10 counter$count = 68607;
	#10 counter$count = 68608;
	#10 counter$count = 68609;
	#10 counter$count = 68610;
	#10 counter$count = 68611;
	#10 counter$count = 68612;
	#10 counter$count = 68613;
	#10 counter$count = 68614;
	#10 counter$count = 68615;
	#10 counter$count = 68616;
	#10 counter$count = 68617;
	#10 counter$count = 68618;
	#10 counter$count = 68619;
	#10 counter$count = 68620;
	#10 counter$count = 68621;
	#10 counter$count = 68622;
	#10 counter$count = 68623;
	#10 counter$count = 68624;
	#10 counter$count = 68625;
	#10 counter$count = 68626;
	#10 counter$count = 68627;
	#10 counter$count = 68628;
	#10 counter$count = 68629;
	#10 counter$count = 68630;
	#10 counter$count = 68631;
	#10 counter$count = 68632;
	#10 counter$count = 68633;
	#10 counter$count = 68634;
	#10 counter$count = 68635;
	#10 counter$count = 68636;
	#10 counter$count = 68637;
	#10 counter$count = 68638;
	#10 counter$count = 68639;
	#10 counter$count = 68640;
	#10 counter$count = 68641;
	#10 counter$count = 68642;
	#10 counter$count = 68643;
	#10 counter$count = 68644;
	#10 counter$count = 68645;
	#10 counter$count = 68646;
	#10 counter$count = 68647;
	#10 counter$count = 68648;
	#10 counter$count = 68649;
	#10 counter$count = 68650;
	#10 counter$count = 68651;
	#10 counter$count = 68652;
	#10 counter$count = 68653;
	#10 counter$count = 68654;
	#10 counter$count = 68655;
	#10 counter$count = 68656;
	#10 counter$count = 68657;
	#10 counter$count = 68658;
	#10 counter$count = 68659;
	#10 counter$count = 68660;
	#10 counter$count = 68661;
	#10 counter$count = 68662;
	#10 counter$count = 68663;
	#10 counter$count = 68664;
	#10 counter$count = 68665;
	#10 counter$count = 68666;
	#10 counter$count = 68667;
	#10 counter$count = 68668;
	#10 counter$count = 68669;
	#10 counter$count = 68670;
	#10 counter$count = 68671;
	#10 counter$count = 68672;
	#10 counter$count = 68673;
	#10 counter$count = 68674;
	#10 counter$count = 68675;
	#10 counter$count = 68676;
	#10 counter$count = 68677;
	#10 counter$count = 68678;
	#10 counter$count = 68679;
	#10 counter$count = 68680;
	#10 counter$count = 68681;
	#10 counter$count = 68682;
	#10 counter$count = 68683;
	#10 counter$count = 68684;
	#10 counter$count = 68685;
	#10 counter$count = 68686;
	#10 counter$count = 68687;
	#10 counter$count = 68688;
	#10 counter$count = 68689;
	#10 counter$count = 68690;
	#10 counter$count = 68691;
	#10 counter$count = 68692;
	#10 counter$count = 68693;
	#10 counter$count = 68694;
	#10 counter$count = 68695;
	#10 counter$count = 68696;
	#10 counter$count = 68697;
	#10 counter$count = 68698;
	#10 counter$count = 68699;
	#10 counter$count = 68700;
	#10 counter$count = 68701;
	#10 counter$count = 68702;
	#10 counter$count = 68703;
	#10 counter$count = 68704;
	#10 counter$count = 68705;
	#10 counter$count = 68706;
	#10 counter$count = 68707;
	#10 counter$count = 68708;
	#10 counter$count = 68709;
	#10 counter$count = 68710;
	#10 counter$count = 68711;
	#10 counter$count = 68712;
	#10 counter$count = 68713;
	#10 counter$count = 68714;
	#10 counter$count = 68715;
	#10 counter$count = 68716;
	#10 counter$count = 68717;
	#10 counter$count = 68718;
	#10 counter$count = 68719;
	#10 counter$count = 68720;
	#10 counter$count = 68721;
	#10 counter$count = 68722;
	#10 counter$count = 68723;
	#10 counter$count = 68724;
	#10 counter$count = 68725;
	#10 counter$count = 68726;
	#10 counter$count = 68727;
	#10 counter$count = 68728;
	#10 counter$count = 68729;
	#10 counter$count = 68730;
	#10 counter$count = 68731;
	#10 counter$count = 68732;
	#10 counter$count = 68733;
	#10 counter$count = 68734;
	#10 counter$count = 68735;
	#10 counter$count = 68736;
	#10 counter$count = 68737;
	#10 counter$count = 68738;
	#10 counter$count = 68739;
	#10 counter$count = 68740;
	#10 counter$count = 68741;
	#10 counter$count = 68742;
	#10 counter$count = 68743;
	#10 counter$count = 68744;
	#10 counter$count = 68745;
	#10 counter$count = 68746;
	#10 counter$count = 68747;
	#10 counter$count = 68748;
	#10 counter$count = 68749;
	#10 counter$count = 68750;
	#10 counter$count = 68751;
	#10 counter$count = 68752;
	#10 counter$count = 68753;
	#10 counter$count = 68754;
	#10 counter$count = 68755;
	#10 counter$count = 68756;
	#10 counter$count = 68757;
	#10 counter$count = 68758;
	#10 counter$count = 68759;
	#10 counter$count = 68760;
	#10 counter$count = 68761;
	#10 counter$count = 68762;
	#10 counter$count = 68763;
	#10 counter$count = 68764;
	#10 counter$count = 68765;
	#10 counter$count = 68766;
	#10 counter$count = 68767;
	#10 counter$count = 68768;
	#10 counter$count = 68769;
	#10 counter$count = 68770;
	#10 counter$count = 68771;
	#10 counter$count = 68772;
	#10 counter$count = 68773;
	#10 counter$count = 68774;
	#10 counter$count = 68775;
	#10 counter$count = 68776;
	#10 counter$count = 68777;
	#10 counter$count = 68778;
	#10 counter$count = 68779;
	#10 counter$count = 68780;
	#10 counter$count = 68781;
	#10 counter$count = 68782;
	#10 counter$count = 68783;
	#10 counter$count = 68784;
	#10 counter$count = 68785;
	#10 counter$count = 68786;
	#10 counter$count = 68787;
	#10 counter$count = 68788;
	#10 counter$count = 68789;
	#10 counter$count = 68790;
	#10 counter$count = 68791;
	#10 counter$count = 68792;
	#10 counter$count = 68793;
	#10 counter$count = 68794;
	#10 counter$count = 68795;
	#10 counter$count = 68796;
	#10 counter$count = 68797;
	#10 counter$count = 68798;
	#10 counter$count = 68799;
	#10 counter$count = 68800;
	#10 counter$count = 68801;
	#10 counter$count = 68802;
	#10 counter$count = 68803;
	#10 counter$count = 68804;
	#10 counter$count = 68805;
	#10 counter$count = 68806;
	#10 counter$count = 68807;
	#10 counter$count = 68808;
	#10 counter$count = 68809;
	#10 counter$count = 68810;
	#10 counter$count = 68811;
	#10 counter$count = 68812;
	#10 counter$count = 68813;
	#10 counter$count = 68814;
	#10 counter$count = 68815;
	#10 counter$count = 68816;
	#10 counter$count = 68817;
	#10 counter$count = 68818;
	#10 counter$count = 68819;
	#10 counter$count = 68820;
	#10 counter$count = 68821;
	#10 counter$count = 68822;
	#10 counter$count = 68823;
	#10 counter$count = 68824;
	#10 counter$count = 68825;
	#10 counter$count = 68826;
	#10 counter$count = 68827;
	#10 counter$count = 68828;
	#10 counter$count = 68829;
	#10 counter$count = 68830;
	#10 counter$count = 68831;
	#10 counter$count = 68832;
	#10 counter$count = 68833;
	#10 counter$count = 68834;
	#10 counter$count = 68835;
	#10 counter$count = 68836;
	#10 counter$count = 68837;
	#10 counter$count = 68838;
	#10 counter$count = 68839;
	#10 counter$count = 68840;
	#10 counter$count = 68841;
	#10 counter$count = 68842;
	#10 counter$count = 68843;
	#10 counter$count = 68844;
	#10 counter$count = 68845;
	#10 counter$count = 68846;
	#10 counter$count = 68847;
	#10 counter$count = 68848;
	#10 counter$count = 68849;
	#10 counter$count = 68850;
	#10 counter$count = 68851;
	#10 counter$count = 68852;
	#10 counter$count = 68853;
	#10 counter$count = 68854;
	#10 counter$count = 68855;
	#10 counter$count = 68856;
	#10 counter$count = 68857;
	#10 counter$count = 68858;
	#10 counter$count = 68859;
	#10 counter$count = 68860;
	#10 counter$count = 68861;
	#10 counter$count = 68862;
	#10 counter$count = 68863;
	#10 counter$count = 68864;
	#10 counter$count = 68865;
	#10 counter$count = 68866;
	#10 counter$count = 68867;
	#10 counter$count = 68868;
	#10 counter$count = 68869;
	#10 counter$count = 68870;
	#10 counter$count = 68871;
	#10 counter$count = 68872;
	#10 counter$count = 68873;
	#10 counter$count = 68874;
	#10 counter$count = 68875;
	#10 counter$count = 68876;
	#10 counter$count = 68877;
	#10 counter$count = 68878;
	#10 counter$count = 68879;
	#10 counter$count = 68880;
	#10 counter$count = 68881;
	#10 counter$count = 68882;
	#10 counter$count = 68883;
	#10 counter$count = 68884;
	#10 counter$count = 68885;
	#10 counter$count = 68886;
	#10 counter$count = 68887;
	#10 counter$count = 68888;
	#10 counter$count = 68889;
	#10 counter$count = 68890;
	#10 counter$count = 68891;
	#10 counter$count = 68892;
	#10 counter$count = 68893;
	#10 counter$count = 68894;
	#10 counter$count = 68895;
	#10 counter$count = 68896;
	#10 counter$count = 68897;
	#10 counter$count = 68898;
	#10 counter$count = 68899;
	#10 counter$count = 68900;
	#10 counter$count = 68901;
	#10 counter$count = 68902;
	#10 counter$count = 68903;
	#10 counter$count = 68904;
	#10 counter$count = 68905;
	#10 counter$count = 68906;
	#10 counter$count = 68907;
	#10 counter$count = 68908;
	#10 counter$count = 68909;
	#10 counter$count = 68910;
	#10 counter$count = 68911;
	#10 counter$count = 68912;
	#10 counter$count = 68913;
	#10 counter$count = 68914;
	#10 counter$count = 68915;
	#10 counter$count = 68916;
	#10 counter$count = 68917;
	#10 counter$count = 68918;
	#10 counter$count = 68919;
	#10 counter$count = 68920;
	#10 counter$count = 68921;
	#10 counter$count = 68922;
	#10 counter$count = 68923;
	#10 counter$count = 68924;
	#10 counter$count = 68925;
	#10 counter$count = 68926;
	#10 counter$count = 68927;
	#10 counter$count = 68928;
	#10 counter$count = 68929;
	#10 counter$count = 68930;
	#10 counter$count = 68931;
	#10 counter$count = 68932;
	#10 counter$count = 68933;
	#10 counter$count = 68934;
	#10 counter$count = 68935;
	#10 counter$count = 68936;
	#10 counter$count = 68937;
	#10 counter$count = 68938;
	#10 counter$count = 68939;
	#10 counter$count = 68940;
	#10 counter$count = 68941;
	#10 counter$count = 68942;
	#10 counter$count = 68943;
	#10 counter$count = 68944;
	#10 counter$count = 68945;
	#10 counter$count = 68946;
	#10 counter$count = 68947;
	#10 counter$count = 68948;
	#10 counter$count = 68949;
	#10 counter$count = 68950;
	#10 counter$count = 68951;
	#10 counter$count = 68952;
	#10 counter$count = 68953;
	#10 counter$count = 68954;
	#10 counter$count = 68955;
	#10 counter$count = 68956;
	#10 counter$count = 68957;
	#10 counter$count = 68958;
	#10 counter$count = 68959;
	#10 counter$count = 68960;
	#10 counter$count = 68961;
	#10 counter$count = 68962;
	#10 counter$count = 68963;
	#10 counter$count = 68964;
	#10 counter$count = 68965;
	#10 counter$count = 68966;
	#10 counter$count = 68967;
	#10 counter$count = 68968;
	#10 counter$count = 68969;
	#10 counter$count = 68970;
	#10 counter$count = 68971;
	#10 counter$count = 68972;
	#10 counter$count = 68973;
	#10 counter$count = 68974;
	#10 counter$count = 68975;
	#10 counter$count = 68976;
	#10 counter$count = 68977;
	#10 counter$count = 68978;
	#10 counter$count = 68979;
	#10 counter$count = 68980;
	#10 counter$count = 68981;
	#10 counter$count = 68982;
	#10 counter$count = 68983;
	#10 counter$count = 68984;
	#10 counter$count = 68985;
	#10 counter$count = 68986;
	#10 counter$count = 68987;
	#10 counter$count = 68988;
	#10 counter$count = 68989;
	#10 counter$count = 68990;
	#10 counter$count = 68991;
	#10 counter$count = 68992;
	#10 counter$count = 68993;
	#10 counter$count = 68994;
	#10 counter$count = 68995;
	#10 counter$count = 68996;
	#10 counter$count = 68997;
	#10 counter$count = 68998;
	#10 counter$count = 68999;
	#10 counter$count = 69000;
	#10 counter$count = 69001;
	#10 counter$count = 69002;
	#10 counter$count = 69003;
	#10 counter$count = 69004;
	#10 counter$count = 69005;
	#10 counter$count = 69006;
	#10 counter$count = 69007;
	#10 counter$count = 69008;
	#10 counter$count = 69009;
	#10 counter$count = 69010;
	#10 counter$count = 69011;
	#10 counter$count = 69012;
	#10 counter$count = 69013;
	#10 counter$count = 69014;
	#10 counter$count = 69015;
	#10 counter$count = 69016;
	#10 counter$count = 69017;
	#10 counter$count = 69018;
	#10 counter$count = 69019;
	#10 counter$count = 69020;
	#10 counter$count = 69021;
	#10 counter$count = 69022;
	#10 counter$count = 69023;
	#10 counter$count = 69024;
	#10 counter$count = 69025;
	#10 counter$count = 69026;
	#10 counter$count = 69027;
	#10 counter$count = 69028;
	#10 counter$count = 69029;
	#10 counter$count = 69030;
	#10 counter$count = 69031;
	#10 counter$count = 69032;
	#10 counter$count = 69033;
	#10 counter$count = 69034;
	#10 counter$count = 69035;
	#10 counter$count = 69036;
	#10 counter$count = 69037;
	#10 counter$count = 69038;
	#10 counter$count = 69039;
	#10 counter$count = 69040;
	#10 counter$count = 69041;
	#10 counter$count = 69042;
	#10 counter$count = 69043;
	#10 counter$count = 69044;
	#10 counter$count = 69045;
	#10 counter$count = 69046;
	#10 counter$count = 69047;
	#10 counter$count = 69048;
	#10 counter$count = 69049;
	#10 counter$count = 69050;
	#10 counter$count = 69051;
	#10 counter$count = 69052;
	#10 counter$count = 69053;
	#10 counter$count = 69054;
	#10 counter$count = 69055;
	#10 counter$count = 69056;
	#10 counter$count = 69057;
	#10 counter$count = 69058;
	#10 counter$count = 69059;
	#10 counter$count = 69060;
	#10 counter$count = 69061;
	#10 counter$count = 69062;
	#10 counter$count = 69063;
	#10 counter$count = 69064;
	#10 counter$count = 69065;
	#10 counter$count = 69066;
	#10 counter$count = 69067;
	#10 counter$count = 69068;
	#10 counter$count = 69069;
	#10 counter$count = 69070;
	#10 counter$count = 69071;
	#10 counter$count = 69072;
	#10 counter$count = 69073;
	#10 counter$count = 69074;
	#10 counter$count = 69075;
	#10 counter$count = 69076;
	#10 counter$count = 69077;
	#10 counter$count = 69078;
	#10 counter$count = 69079;
	#10 counter$count = 69080;
	#10 counter$count = 69081;
	#10 counter$count = 69082;
	#10 counter$count = 69083;
	#10 counter$count = 69084;
	#10 counter$count = 69085;
	#10 counter$count = 69086;
	#10 counter$count = 69087;
	#10 counter$count = 69088;
	#10 counter$count = 69089;
	#10 counter$count = 69090;
	#10 counter$count = 69091;
	#10 counter$count = 69092;
	#10 counter$count = 69093;
	#10 counter$count = 69094;
	#10 counter$count = 69095;
	#10 counter$count = 69096;
	#10 counter$count = 69097;
	#10 counter$count = 69098;
	#10 counter$count = 69099;
	#10 counter$count = 69100;
	#10 counter$count = 69101;
	#10 counter$count = 69102;
	#10 counter$count = 69103;
	#10 counter$count = 69104;
	#10 counter$count = 69105;
	#10 counter$count = 69106;
	#10 counter$count = 69107;
	#10 counter$count = 69108;
	#10 counter$count = 69109;
	#10 counter$count = 69110;
	#10 counter$count = 69111;
	#10 counter$count = 69112;
	#10 counter$count = 69113;
	#10 counter$count = 69114;
	#10 counter$count = 69115;
	#10 counter$count = 69116;
	#10 counter$count = 69117;
	#10 counter$count = 69118;
	#10 counter$count = 69119;
	#10 counter$count = 69120;
	#10 counter$count = 69121;
	#10 counter$count = 69122;
	#10 counter$count = 69123;
	#10 counter$count = 69124;
	#10 counter$count = 69125;
	#10 counter$count = 69126;
	#10 counter$count = 69127;
	#10 counter$count = 69128;
	#10 counter$count = 69129;
	#10 counter$count = 69130;
	#10 counter$count = 69131;
	#10 counter$count = 69132;
	#10 counter$count = 69133;
	#10 counter$count = 69134;
	#10 counter$count = 69135;
	#10 counter$count = 69136;
	#10 counter$count = 69137;
	#10 counter$count = 69138;
	#10 counter$count = 69139;
	#10 counter$count = 69140;
	#10 counter$count = 69141;
	#10 counter$count = 69142;
	#10 counter$count = 69143;
	#10 counter$count = 69144;
	#10 counter$count = 69145;
	#10 counter$count = 69146;
	#10 counter$count = 69147;
	#10 counter$count = 69148;
	#10 counter$count = 69149;
	#10 counter$count = 69150;
	#10 counter$count = 69151;
	#10 counter$count = 69152;
	#10 counter$count = 69153;
	#10 counter$count = 69154;
	#10 counter$count = 69155;
	#10 counter$count = 69156;
	#10 counter$count = 69157;
	#10 counter$count = 69158;
	#10 counter$count = 69159;
	#10 counter$count = 69160;
	#10 counter$count = 69161;
	#10 counter$count = 69162;
	#10 counter$count = 69163;
	#10 counter$count = 69164;
	#10 counter$count = 69165;
	#10 counter$count = 69166;
	#10 counter$count = 69167;
	#10 counter$count = 69168;
	#10 counter$count = 69169;
	#10 counter$count = 69170;
	#10 counter$count = 69171;
	#10 counter$count = 69172;
	#10 counter$count = 69173;
	#10 counter$count = 69174;
	#10 counter$count = 69175;
	#10 counter$count = 69176;
	#10 counter$count = 69177;
	#10 counter$count = 69178;
	#10 counter$count = 69179;
	#10 counter$count = 69180;
	#10 counter$count = 69181;
	#10 counter$count = 69182;
	#10 counter$count = 69183;
	#10 counter$count = 69184;
	#10 counter$count = 69185;
	#10 counter$count = 69186;
	#10 counter$count = 69187;
	#10 counter$count = 69188;
	#10 counter$count = 69189;
	#10 counter$count = 69190;
	#10 counter$count = 69191;
	#10 counter$count = 69192;
	#10 counter$count = 69193;
	#10 counter$count = 69194;
	#10 counter$count = 69195;
	#10 counter$count = 69196;
	#10 counter$count = 69197;
	#10 counter$count = 69198;
	#10 counter$count = 69199;
	#10 counter$count = 69200;
	#10 counter$count = 69201;
	#10 counter$count = 69202;
	#10 counter$count = 69203;
	#10 counter$count = 69204;
	#10 counter$count = 69205;
	#10 counter$count = 69206;
	#10 counter$count = 69207;
	#10 counter$count = 69208;
	#10 counter$count = 69209;
	#10 counter$count = 69210;
	#10 counter$count = 69211;
	#10 counter$count = 69212;
	#10 counter$count = 69213;
	#10 counter$count = 69214;
	#10 counter$count = 69215;
	#10 counter$count = 69216;
	#10 counter$count = 69217;
	#10 counter$count = 69218;
	#10 counter$count = 69219;
	#10 counter$count = 69220;
	#10 counter$count = 69221;
	#10 counter$count = 69222;
	#10 counter$count = 69223;
	#10 counter$count = 69224;
	#10 counter$count = 69225;
	#10 counter$count = 69226;
	#10 counter$count = 69227;
	#10 counter$count = 69228;
	#10 counter$count = 69229;
	#10 counter$count = 69230;
	#10 counter$count = 69231;
	#10 counter$count = 69232;
	#10 counter$count = 69233;
	#10 counter$count = 69234;
	#10 counter$count = 69235;
	#10 counter$count = 69236;
	#10 counter$count = 69237;
	#10 counter$count = 69238;
	#10 counter$count = 69239;
	#10 counter$count = 69240;
	#10 counter$count = 69241;
	#10 counter$count = 69242;
	#10 counter$count = 69243;
	#10 counter$count = 69244;
	#10 counter$count = 69245;
	#10 counter$count = 69246;
	#10 counter$count = 69247;
	#10 counter$count = 69248;
	#10 counter$count = 69249;
	#10 counter$count = 69250;
	#10 counter$count = 69251;
	#10 counter$count = 69252;
	#10 counter$count = 69253;
	#10 counter$count = 69254;
	#10 counter$count = 69255;
	#10 counter$count = 69256;
	#10 counter$count = 69257;
	#10 counter$count = 69258;
	#10 counter$count = 69259;
	#10 counter$count = 69260;
	#10 counter$count = 69261;
	#10 counter$count = 69262;
	#10 counter$count = 69263;
	#10 counter$count = 69264;
	#10 counter$count = 69265;
	#10 counter$count = 69266;
	#10 counter$count = 69267;
	#10 counter$count = 69268;
	#10 counter$count = 69269;
	#10 counter$count = 69270;
	#10 counter$count = 69271;
	#10 counter$count = 69272;
	#10 counter$count = 69273;
	#10 counter$count = 69274;
	#10 counter$count = 69275;
	#10 counter$count = 69276;
	#10 counter$count = 69277;
	#10 counter$count = 69278;
	#10 counter$count = 69279;
	#10 counter$count = 69280;
	#10 counter$count = 69281;
	#10 counter$count = 69282;
	#10 counter$count = 69283;
	#10 counter$count = 69284;
	#10 counter$count = 69285;
	#10 counter$count = 69286;
	#10 counter$count = 69287;
	#10 counter$count = 69288;
	#10 counter$count = 69289;
	#10 counter$count = 69290;
	#10 counter$count = 69291;
	#10 counter$count = 69292;
	#10 counter$count = 69293;
	#10 counter$count = 69294;
	#10 counter$count = 69295;
	#10 counter$count = 69296;
	#10 counter$count = 69297;
	#10 counter$count = 69298;
	#10 counter$count = 69299;
	#10 counter$count = 69300;
	#10 counter$count = 69301;
	#10 counter$count = 69302;
	#10 counter$count = 69303;
	#10 counter$count = 69304;
	#10 counter$count = 69305;
	#10 counter$count = 69306;
	#10 counter$count = 69307;
	#10 counter$count = 69308;
	#10 counter$count = 69309;
	#10 counter$count = 69310;
	#10 counter$count = 69311;
	#10 counter$count = 69312;
	#10 counter$count = 69313;
	#10 counter$count = 69314;
	#10 counter$count = 69315;
	#10 counter$count = 69316;
	#10 counter$count = 69317;
	#10 counter$count = 69318;
	#10 counter$count = 69319;
	#10 counter$count = 69320;
	#10 counter$count = 69321;
	#10 counter$count = 69322;
	#10 counter$count = 69323;
	#10 counter$count = 69324;
	#10 counter$count = 69325;
	#10 counter$count = 69326;
	#10 counter$count = 69327;
	#10 counter$count = 69328;
	#10 counter$count = 69329;
	#10 counter$count = 69330;
	#10 counter$count = 69331;
	#10 counter$count = 69332;
	#10 counter$count = 69333;
	#10 counter$count = 69334;
	#10 counter$count = 69335;
	#10 counter$count = 69336;
	#10 counter$count = 69337;
	#10 counter$count = 69338;
	#10 counter$count = 69339;
	#10 counter$count = 69340;
	#10 counter$count = 69341;
	#10 counter$count = 69342;
	#10 counter$count = 69343;
	#10 counter$count = 69344;
	#10 counter$count = 69345;
	#10 counter$count = 69346;
	#10 counter$count = 69347;
	#10 counter$count = 69348;
	#10 counter$count = 69349;
	#10 counter$count = 69350;
	#10 counter$count = 69351;
	#10 counter$count = 69352;
	#10 counter$count = 69353;
	#10 counter$count = 69354;
	#10 counter$count = 69355;
	#10 counter$count = 69356;
	#10 counter$count = 69357;
	#10 counter$count = 69358;
	#10 counter$count = 69359;
	#10 counter$count = 69360;
	#10 counter$count = 69361;
	#10 counter$count = 69362;
	#10 counter$count = 69363;
	#10 counter$count = 69364;
	#10 counter$count = 69365;
	#10 counter$count = 69366;
	#10 counter$count = 69367;
	#10 counter$count = 69368;
	#10 counter$count = 69369;
	#10 counter$count = 69370;
	#10 counter$count = 69371;
	#10 counter$count = 69372;
	#10 counter$count = 69373;
	#10 counter$count = 69374;
	#10 counter$count = 69375;
	#10 counter$count = 69376;
	#10 counter$count = 69377;
	#10 counter$count = 69378;
	#10 counter$count = 69379;
	#10 counter$count = 69380;
	#10 counter$count = 69381;
	#10 counter$count = 69382;
	#10 counter$count = 69383;
	#10 counter$count = 69384;
	#10 counter$count = 69385;
	#10 counter$count = 69386;
	#10 counter$count = 69387;
	#10 counter$count = 69388;
	#10 counter$count = 69389;
	#10 counter$count = 69390;
	#10 counter$count = 69391;
	#10 counter$count = 69392;
	#10 counter$count = 69393;
	#10 counter$count = 69394;
	#10 counter$count = 69395;
	#10 counter$count = 69396;
	#10 counter$count = 69397;
	#10 counter$count = 69398;
	#10 counter$count = 69399;
	#10 counter$count = 69400;
	#10 counter$count = 69401;
	#10 counter$count = 69402;
	#10 counter$count = 69403;
	#10 counter$count = 69404;
	#10 counter$count = 69405;
	#10 counter$count = 69406;
	#10 counter$count = 69407;
	#10 counter$count = 69408;
	#10 counter$count = 69409;
	#10 counter$count = 69410;
	#10 counter$count = 69411;
	#10 counter$count = 69412;
	#10 counter$count = 69413;
	#10 counter$count = 69414;
	#10 counter$count = 69415;
	#10 counter$count = 69416;
	#10 counter$count = 69417;
	#10 counter$count = 69418;
	#10 counter$count = 69419;
	#10 counter$count = 69420;
	#10 counter$count = 69421;
	#10 counter$count = 69422;
	#10 counter$count = 69423;
	#10 counter$count = 69424;
	#10 counter$count = 69425;
	#10 counter$count = 69426;
	#10 counter$count = 69427;
	#10 counter$count = 69428;
	#10 counter$count = 69429;
	#10 counter$count = 69430;
	#10 counter$count = 69431;
	#10 counter$count = 69432;
	#10 counter$count = 69433;
	#10 counter$count = 69434;
	#10 counter$count = 69435;
	#10 counter$count = 69436;
	#10 counter$count = 69437;
	#10 counter$count = 69438;
	#10 counter$count = 69439;
	#10 counter$count = 69440;
	#10 counter$count = 69441;
	#10 counter$count = 69442;
	#10 counter$count = 69443;
	#10 counter$count = 69444;
	#10 counter$count = 69445;
	#10 counter$count = 69446;
	#10 counter$count = 69447;
	#10 counter$count = 69448;
	#10 counter$count = 69449;
	#10 counter$count = 69450;
	#10 counter$count = 69451;
	#10 counter$count = 69452;
	#10 counter$count = 69453;
	#10 counter$count = 69454;
	#10 counter$count = 69455;
	#10 counter$count = 69456;
	#10 counter$count = 69457;
	#10 counter$count = 69458;
	#10 counter$count = 69459;
	#10 counter$count = 69460;
	#10 counter$count = 69461;
	#10 counter$count = 69462;
	#10 counter$count = 69463;
	#10 counter$count = 69464;
	#10 counter$count = 69465;
	#10 counter$count = 69466;
	#10 counter$count = 69467;
	#10 counter$count = 69468;
	#10 counter$count = 69469;
	#10 counter$count = 69470;
	#10 counter$count = 69471;
	#10 counter$count = 69472;
	#10 counter$count = 69473;
	#10 counter$count = 69474;
	#10 counter$count = 69475;
	#10 counter$count = 69476;
	#10 counter$count = 69477;
	#10 counter$count = 69478;
	#10 counter$count = 69479;
	#10 counter$count = 69480;
	#10 counter$count = 69481;
	#10 counter$count = 69482;
	#10 counter$count = 69483;
	#10 counter$count = 69484;
	#10 counter$count = 69485;
	#10 counter$count = 69486;
	#10 counter$count = 69487;
	#10 counter$count = 69488;
	#10 counter$count = 69489;
	#10 counter$count = 69490;
	#10 counter$count = 69491;
	#10 counter$count = 69492;
	#10 counter$count = 69493;
	#10 counter$count = 69494;
	#10 counter$count = 69495;
	#10 counter$count = 69496;
	#10 counter$count = 69497;
	#10 counter$count = 69498;
	#10 counter$count = 69499;
	#10 counter$count = 69500;
	#10 counter$count = 69501;
	#10 counter$count = 69502;
	#10 counter$count = 69503;
	#10 counter$count = 69504;
	#10 counter$count = 69505;
	#10 counter$count = 69506;
	#10 counter$count = 69507;
	#10 counter$count = 69508;
	#10 counter$count = 69509;
	#10 counter$count = 69510;
	#10 counter$count = 69511;
	#10 counter$count = 69512;
	#10 counter$count = 69513;
	#10 counter$count = 69514;
	#10 counter$count = 69515;
	#10 counter$count = 69516;
	#10 counter$count = 69517;
	#10 counter$count = 69518;
	#10 counter$count = 69519;
	#10 counter$count = 69520;
	#10 counter$count = 69521;
	#10 counter$count = 69522;
	#10 counter$count = 69523;
	#10 counter$count = 69524;
	#10 counter$count = 69525;
	#10 counter$count = 69526;
	#10 counter$count = 69527;
	#10 counter$count = 69528;
	#10 counter$count = 69529;
	#10 counter$count = 69530;
	#10 counter$count = 69531;
	#10 counter$count = 69532;
	#10 counter$count = 69533;
	#10 counter$count = 69534;
	#10 counter$count = 69535;
	#10 counter$count = 69536;
	#10 counter$count = 69537;
	#10 counter$count = 69538;
	#10 counter$count = 69539;
	#10 counter$count = 69540;
	#10 counter$count = 69541;
	#10 counter$count = 69542;
	#10 counter$count = 69543;
	#10 counter$count = 69544;
	#10 counter$count = 69545;
	#10 counter$count = 69546;
	#10 counter$count = 69547;
	#10 counter$count = 69548;
	#10 counter$count = 69549;
	#10 counter$count = 69550;
	#10 counter$count = 69551;
	#10 counter$count = 69552;
	#10 counter$count = 69553;
	#10 counter$count = 69554;
	#10 counter$count = 69555;
	#10 counter$count = 69556;
	#10 counter$count = 69557;
	#10 counter$count = 69558;
	#10 counter$count = 69559;
	#10 counter$count = 69560;
	#10 counter$count = 69561;
	#10 counter$count = 69562;
	#10 counter$count = 69563;
	#10 counter$count = 69564;
	#10 counter$count = 69565;
	#10 counter$count = 69566;
	#10 counter$count = 69567;
	#10 counter$count = 69568;
	#10 counter$count = 69569;
	#10 counter$count = 69570;
	#10 counter$count = 69571;
	#10 counter$count = 69572;
	#10 counter$count = 69573;
	#10 counter$count = 69574;
	#10 counter$count = 69575;
	#10 counter$count = 69576;
	#10 counter$count = 69577;
	#10 counter$count = 69578;
	#10 counter$count = 69579;
	#10 counter$count = 69580;
	#10 counter$count = 69581;
	#10 counter$count = 69582;
	#10 counter$count = 69583;
	#10 counter$count = 69584;
	#10 counter$count = 69585;
	#10 counter$count = 69586;
	#10 counter$count = 69587;
	#10 counter$count = 69588;
	#10 counter$count = 69589;
	#10 counter$count = 69590;
	#10 counter$count = 69591;
	#10 counter$count = 69592;
	#10 counter$count = 69593;
	#10 counter$count = 69594;
	#10 counter$count = 69595;
	#10 counter$count = 69596;
	#10 counter$count = 69597;
	#10 counter$count = 69598;
	#10 counter$count = 69599;
	#10 counter$count = 69600;
	#10 counter$count = 69601;
	#10 counter$count = 69602;
	#10 counter$count = 69603;
	#10 counter$count = 69604;
	#10 counter$count = 69605;
	#10 counter$count = 69606;
	#10 counter$count = 69607;
	#10 counter$count = 69608;
	#10 counter$count = 69609;
	#10 counter$count = 69610;
	#10 counter$count = 69611;
	#10 counter$count = 69612;
	#10 counter$count = 69613;
	#10 counter$count = 69614;
	#10 counter$count = 69615;
	#10 counter$count = 69616;
	#10 counter$count = 69617;
	#10 counter$count = 69618;
	#10 counter$count = 69619;
	#10 counter$count = 69620;
	#10 counter$count = 69621;
	#10 counter$count = 69622;
	#10 counter$count = 69623;
	#10 counter$count = 69624;
	#10 counter$count = 69625;
	#10 counter$count = 69626;
	#10 counter$count = 69627;
	#10 counter$count = 69628;
	#10 counter$count = 69629;
	#10 counter$count = 69630;
	#10 counter$count = 69631;
	#10 counter$count = 69632;
	#10 counter$count = 69633;
	#10 counter$count = 69634;
	#10 counter$count = 69635;
	#10 counter$count = 69636;
	#10 counter$count = 69637;
	#10 counter$count = 69638;
	#10 counter$count = 69639;
	#10 counter$count = 69640;
	#10 counter$count = 69641;
	#10 counter$count = 69642;
	#10 counter$count = 69643;
	#10 counter$count = 69644;
	#10 counter$count = 69645;
	#10 counter$count = 69646;
	#10 counter$count = 69647;
	#10 counter$count = 69648;
	#10 counter$count = 69649;
	#10 counter$count = 69650;
	#10 counter$count = 69651;
	#10 counter$count = 69652;
	#10 counter$count = 69653;
	#10 counter$count = 69654;
	#10 counter$count = 69655;
	#10 counter$count = 69656;
	#10 counter$count = 69657;
	#10 counter$count = 69658;
	#10 counter$count = 69659;
	#10 counter$count = 69660;
	#10 counter$count = 69661;
	#10 counter$count = 69662;
	#10 counter$count = 69663;
	#10 counter$count = 69664;
	#10 counter$count = 69665;
	#10 counter$count = 69666;
	#10 counter$count = 69667;
	#10 counter$count = 69668;
	#10 counter$count = 69669;
	#10 counter$count = 69670;
	#10 counter$count = 69671;
	#10 counter$count = 69672;
	#10 counter$count = 69673;
	#10 counter$count = 69674;
	#10 counter$count = 69675;
	#10 counter$count = 69676;
	#10 counter$count = 69677;
	#10 counter$count = 69678;
	#10 counter$count = 69679;
	#10 counter$count = 69680;
	#10 counter$count = 69681;
	#10 counter$count = 69682;
	#10 counter$count = 69683;
	#10 counter$count = 69684;
	#10 counter$count = 69685;
	#10 counter$count = 69686;
	#10 counter$count = 69687;
	#10 counter$count = 69688;
	#10 counter$count = 69689;
	#10 counter$count = 69690;
	#10 counter$count = 69691;
	#10 counter$count = 69692;
	#10 counter$count = 69693;
	#10 counter$count = 69694;
	#10 counter$count = 69695;
	#10 counter$count = 69696;
	#10 counter$count = 69697;
	#10 counter$count = 69698;
	#10 counter$count = 69699;
	#10 counter$count = 69700;
	#10 counter$count = 69701;
	#10 counter$count = 69702;
	#10 counter$count = 69703;
	#10 counter$count = 69704;
	#10 counter$count = 69705;
	#10 counter$count = 69706;
	#10 counter$count = 69707;
	#10 counter$count = 69708;
	#10 counter$count = 69709;
	#10 counter$count = 69710;
	#10 counter$count = 69711;
	#10 counter$count = 69712;
	#10 counter$count = 69713;
	#10 counter$count = 69714;
	#10 counter$count = 69715;
	#10 counter$count = 69716;
	#10 counter$count = 69717;
	#10 counter$count = 69718;
	#10 counter$count = 69719;
	#10 counter$count = 69720;
	#10 counter$count = 69721;
	#10 counter$count = 69722;
	#10 counter$count = 69723;
	#10 counter$count = 69724;
	#10 counter$count = 69725;
	#10 counter$count = 69726;
	#10 counter$count = 69727;
	#10 counter$count = 69728;
	#10 counter$count = 69729;
	#10 counter$count = 69730;
	#10 counter$count = 69731;
	#10 counter$count = 69732;
	#10 counter$count = 69733;
	#10 counter$count = 69734;
	#10 counter$count = 69735;
	#10 counter$count = 69736;
	#10 counter$count = 69737;
	#10 counter$count = 69738;
	#10 counter$count = 69739;
	#10 counter$count = 69740;
	#10 counter$count = 69741;
	#10 counter$count = 69742;
	#10 counter$count = 69743;
	#10 counter$count = 69744;
	#10 counter$count = 69745;
	#10 counter$count = 69746;
	#10 counter$count = 69747;
	#10 counter$count = 69748;
	#10 counter$count = 69749;
	#10 counter$count = 69750;
	#10 counter$count = 69751;
	#10 counter$count = 69752;
	#10 counter$count = 69753;
	#10 counter$count = 69754;
	#10 counter$count = 69755;
	#10 counter$count = 69756;
	#10 counter$count = 69757;
	#10 counter$count = 69758;
	#10 counter$count = 69759;
	#10 counter$count = 69760;
	#10 counter$count = 69761;
	#10 counter$count = 69762;
	#10 counter$count = 69763;
	#10 counter$count = 69764;
	#10 counter$count = 69765;
	#10 counter$count = 69766;
	#10 counter$count = 69767;
	#10 counter$count = 69768;
	#10 counter$count = 69769;
	#10 counter$count = 69770;
	#10 counter$count = 69771;
	#10 counter$count = 69772;
	#10 counter$count = 69773;
	#10 counter$count = 69774;
	#10 counter$count = 69775;
	#10 counter$count = 69776;
	#10 counter$count = 69777;
	#10 counter$count = 69778;
	#10 counter$count = 69779;
	#10 counter$count = 69780;
	#10 counter$count = 69781;
	#10 counter$count = 69782;
	#10 counter$count = 69783;
	#10 counter$count = 69784;
	#10 counter$count = 69785;
	#10 counter$count = 69786;
	#10 counter$count = 69787;
	#10 counter$count = 69788;
	#10 counter$count = 69789;
	#10 counter$count = 69790;
	#10 counter$count = 69791;
	#10 counter$count = 69792;
	#10 counter$count = 69793;
	#10 counter$count = 69794;
	#10 counter$count = 69795;
	#10 counter$count = 69796;
	#10 counter$count = 69797;
	#10 counter$count = 69798;
	#10 counter$count = 69799;
	#10 counter$count = 69800;
	#10 counter$count = 69801;
	#10 counter$count = 69802;
	#10 counter$count = 69803;
	#10 counter$count = 69804;
	#10 counter$count = 69805;
	#10 counter$count = 69806;
	#10 counter$count = 69807;
	#10 counter$count = 69808;
	#10 counter$count = 69809;
	#10 counter$count = 69810;
	#10 counter$count = 69811;
	#10 counter$count = 69812;
	#10 counter$count = 69813;
	#10 counter$count = 69814;
	#10 counter$count = 69815;
	#10 counter$count = 69816;
	#10 counter$count = 69817;
	#10 counter$count = 69818;
	#10 counter$count = 69819;
	#10 counter$count = 69820;
	#10 counter$count = 69821;
	#10 counter$count = 69822;
	#10 counter$count = 69823;
	#10 counter$count = 69824;
	#10 counter$count = 69825;
	#10 counter$count = 69826;
	#10 counter$count = 69827;
	#10 counter$count = 69828;
	#10 counter$count = 69829;
	#10 counter$count = 69830;
	#10 counter$count = 69831;
	#10 counter$count = 69832;
	#10 counter$count = 69833;
	#10 counter$count = 69834;
	#10 counter$count = 69835;
	#10 counter$count = 69836;
	#10 counter$count = 69837;
	#10 counter$count = 69838;
	#10 counter$count = 69839;
	#10 counter$count = 69840;
	#10 counter$count = 69841;
	#10 counter$count = 69842;
	#10 counter$count = 69843;
	#10 counter$count = 69844;
	#10 counter$count = 69845;
	#10 counter$count = 69846;
	#10 counter$count = 69847;
	#10 counter$count = 69848;
	#10 counter$count = 69849;
	#10 counter$count = 69850;
	#10 counter$count = 69851;
	#10 counter$count = 69852;
	#10 counter$count = 69853;
	#10 counter$count = 69854;
	#10 counter$count = 69855;
	#10 counter$count = 69856;
	#10 counter$count = 69857;
	#10 counter$count = 69858;
	#10 counter$count = 69859;
	#10 counter$count = 69860;
	#10 counter$count = 69861;
	#10 counter$count = 69862;
	#10 counter$count = 69863;
	#10 counter$count = 69864;
	#10 counter$count = 69865;
	#10 counter$count = 69866;
	#10 counter$count = 69867;
	#10 counter$count = 69868;
	#10 counter$count = 69869;
	#10 counter$count = 69870;
	#10 counter$count = 69871;
	#10 counter$count = 69872;
	#10 counter$count = 69873;
	#10 counter$count = 69874;
	#10 counter$count = 69875;
	#10 counter$count = 69876;
	#10 counter$count = 69877;
	#10 counter$count = 69878;
	#10 counter$count = 69879;
	#10 counter$count = 69880;
	#10 counter$count = 69881;
	#10 counter$count = 69882;
	#10 counter$count = 69883;
	#10 counter$count = 69884;
	#10 counter$count = 69885;
	#10 counter$count = 69886;
	#10 counter$count = 69887;
	#10 counter$count = 69888;
	#10 counter$count = 69889;
	#10 counter$count = 69890;
	#10 counter$count = 69891;
	#10 counter$count = 69892;
	#10 counter$count = 69893;
	#10 counter$count = 69894;
	#10 counter$count = 69895;
	#10 counter$count = 69896;
	#10 counter$count = 69897;
	#10 counter$count = 69898;
	#10 counter$count = 69899;
	#10 counter$count = 69900;
	#10 counter$count = 69901;
	#10 counter$count = 69902;
	#10 counter$count = 69903;
	#10 counter$count = 69904;
	#10 counter$count = 69905;
	#10 counter$count = 69906;
	#10 counter$count = 69907;
	#10 counter$count = 69908;
	#10 counter$count = 69909;
	#10 counter$count = 69910;
	#10 counter$count = 69911;
	#10 counter$count = 69912;
	#10 counter$count = 69913;
	#10 counter$count = 69914;
	#10 counter$count = 69915;
	#10 counter$count = 69916;
	#10 counter$count = 69917;
	#10 counter$count = 69918;
	#10 counter$count = 69919;
	#10 counter$count = 69920;
	#10 counter$count = 69921;
	#10 counter$count = 69922;
	#10 counter$count = 69923;
	#10 counter$count = 69924;
	#10 counter$count = 69925;
	#10 counter$count = 69926;
	#10 counter$count = 69927;
	#10 counter$count = 69928;
	#10 counter$count = 69929;
	#10 counter$count = 69930;
	#10 counter$count = 69931;
	#10 counter$count = 69932;
	#10 counter$count = 69933;
	#10 counter$count = 69934;
	#10 counter$count = 69935;
	#10 counter$count = 69936;
	#10 counter$count = 69937;
	#10 counter$count = 69938;
	#10 counter$count = 69939;
	#10 counter$count = 69940;
	#10 counter$count = 69941;
	#10 counter$count = 69942;
	#10 counter$count = 69943;
	#10 counter$count = 69944;
	#10 counter$count = 69945;
	#10 counter$count = 69946;
	#10 counter$count = 69947;
	#10 counter$count = 69948;
	#10 counter$count = 69949;
	#10 counter$count = 69950;
	#10 counter$count = 69951;
	#10 counter$count = 69952;
	#10 counter$count = 69953;
	#10 counter$count = 69954;
	#10 counter$count = 69955;
	#10 counter$count = 69956;
	#10 counter$count = 69957;
	#10 counter$count = 69958;
	#10 counter$count = 69959;
	#10 counter$count = 69960;
	#10 counter$count = 69961;
	#10 counter$count = 69962;
	#10 counter$count = 69963;
	#10 counter$count = 69964;
	#10 counter$count = 69965;
	#10 counter$count = 69966;
	#10 counter$count = 69967;
	#10 counter$count = 69968;
	#10 counter$count = 69969;
	#10 counter$count = 69970;
	#10 counter$count = 69971;
	#10 counter$count = 69972;
	#10 counter$count = 69973;
	#10 counter$count = 69974;
	#10 counter$count = 69975;
	#10 counter$count = 69976;
	#10 counter$count = 69977;
	#10 counter$count = 69978;
	#10 counter$count = 69979;
	#10 counter$count = 69980;
	#10 counter$count = 69981;
	#10 counter$count = 69982;
	#10 counter$count = 69983;
	#10 counter$count = 69984;
	#10 counter$count = 69985;
	#10 counter$count = 69986;
	#10 counter$count = 69987;
	#10 counter$count = 69988;
	#10 counter$count = 69989;
	#10 counter$count = 69990;
	#10 counter$count = 69991;
	#10 counter$count = 69992;
	#10 counter$count = 69993;
	#10 counter$count = 69994;
	#10 counter$count = 69995;
	#10 counter$count = 69996;
	#10 counter$count = 69997;
	#10 counter$count = 69998;
	#10 counter$count = 69999;
	#10 counter$count = 70000;
	#10 counter$count = 70001;
	#10 counter$count = 70002;
	#10 counter$count = 70003;
	#10 counter$count = 70004;
	#10 counter$count = 70005;
	#10 counter$count = 70006;
	#10 counter$count = 70007;
	#10 counter$count = 70008;
	#10 counter$count = 70009;
	#10 counter$count = 70010;
	#10 counter$count = 70011;
	#10 counter$count = 70012;
	#10 counter$count = 70013;
	#10 counter$count = 70014;
	#10 counter$count = 70015;
	#10 counter$count = 70016;
	#10 counter$count = 70017;
	#10 counter$count = 70018;
	#10 counter$count = 70019;
	#10 counter$count = 70020;
	#10 counter$count = 70021;
	#10 counter$count = 70022;
	#10 counter$count = 70023;
	#10 counter$count = 70024;
	#10 counter$count = 70025;
	#10 counter$count = 70026;
	#10 counter$count = 70027;
	#10 counter$count = 70028;
	#10 counter$count = 70029;
	#10 counter$count = 70030;
	#10 counter$count = 70031;
	#10 counter$count = 70032;
	#10 counter$count = 70033;
	#10 counter$count = 70034;
	#10 counter$count = 70035;
	#10 counter$count = 70036;
	#10 counter$count = 70037;
	#10 counter$count = 70038;
	#10 counter$count = 70039;
	#10 counter$count = 70040;
	#10 counter$count = 70041;
	#10 counter$count = 70042;
	#10 counter$count = 70043;
	#10 counter$count = 70044;
	#10 counter$count = 70045;
	#10 counter$count = 70046;
	#10 counter$count = 70047;
	#10 counter$count = 70048;
	#10 counter$count = 70049;
	#10 counter$count = 70050;
	#10 counter$count = 70051;
	#10 counter$count = 70052;
	#10 counter$count = 70053;
	#10 counter$count = 70054;
	#10 counter$count = 70055;
	#10 counter$count = 70056;
	#10 counter$count = 70057;
	#10 counter$count = 70058;
	#10 counter$count = 70059;
	#10 counter$count = 70060;
	#10 counter$count = 70061;
	#10 counter$count = 70062;
	#10 counter$count = 70063;
	#10 counter$count = 70064;
	#10 counter$count = 70065;
	#10 counter$count = 70066;
	#10 counter$count = 70067;
	#10 counter$count = 70068;
	#10 counter$count = 70069;
	#10 counter$count = 70070;
	#10 counter$count = 70071;
	#10 counter$count = 70072;
	#10 counter$count = 70073;
	#10 counter$count = 70074;
	#10 counter$count = 70075;
	#10 counter$count = 70076;
	#10 counter$count = 70077;
	#10 counter$count = 70078;
	#10 counter$count = 70079;
	#10 counter$count = 70080;
	#10 counter$count = 70081;
	#10 counter$count = 70082;
	#10 counter$count = 70083;
	#10 counter$count = 70084;
	#10 counter$count = 70085;
	#10 counter$count = 70086;
	#10 counter$count = 70087;
	#10 counter$count = 70088;
	#10 counter$count = 70089;
	#10 counter$count = 70090;
	#10 counter$count = 70091;
	#10 counter$count = 70092;
	#10 counter$count = 70093;
	#10 counter$count = 70094;
	#10 counter$count = 70095;
	#10 counter$count = 70096;
	#10 counter$count = 70097;
	#10 counter$count = 70098;
	#10 counter$count = 70099;
	#10 counter$count = 70100;
	#10 counter$count = 70101;
	#10 counter$count = 70102;
	#10 counter$count = 70103;
	#10 counter$count = 70104;
	#10 counter$count = 70105;
	#10 counter$count = 70106;
	#10 counter$count = 70107;
	#10 counter$count = 70108;
	#10 counter$count = 70109;
	#10 counter$count = 70110;
	#10 counter$count = 70111;
	#10 counter$count = 70112;
	#10 counter$count = 70113;
	#10 counter$count = 70114;
	#10 counter$count = 70115;
	#10 counter$count = 70116;
	#10 counter$count = 70117;
	#10 counter$count = 70118;
	#10 counter$count = 70119;
	#10 counter$count = 70120;
	#10 counter$count = 70121;
	#10 counter$count = 70122;
	#10 counter$count = 70123;
	#10 counter$count = 70124;
	#10 counter$count = 70125;
	#10 counter$count = 70126;
	#10 counter$count = 70127;
	#10 counter$count = 70128;
	#10 counter$count = 70129;
	#10 counter$count = 70130;
	#10 counter$count = 70131;
	#10 counter$count = 70132;
	#10 counter$count = 70133;
	#10 counter$count = 70134;
	#10 counter$count = 70135;
	#10 counter$count = 70136;
	#10 counter$count = 70137;
	#10 counter$count = 70138;
	#10 counter$count = 70139;
	#10 counter$count = 70140;
	#10 counter$count = 70141;
	#10 counter$count = 70142;
	#10 counter$count = 70143;
	#10 counter$count = 70144;
	#10 counter$count = 70145;
	#10 counter$count = 70146;
	#10 counter$count = 70147;
	#10 counter$count = 70148;
	#10 counter$count = 70149;
	#10 counter$count = 70150;
	#10 counter$count = 70151;
	#10 counter$count = 70152;
	#10 counter$count = 70153;
	#10 counter$count = 70154;
	#10 counter$count = 70155;
	#10 counter$count = 70156;
	#10 counter$count = 70157;
	#10 counter$count = 70158;
	#10 counter$count = 70159;
	#10 counter$count = 70160;
	#10 counter$count = 70161;
	#10 counter$count = 70162;
	#10 counter$count = 70163;
	#10 counter$count = 70164;
	#10 counter$count = 70165;
	#10 counter$count = 70166;
	#10 counter$count = 70167;
	#10 counter$count = 70168;
	#10 counter$count = 70169;
	#10 counter$count = 70170;
	#10 counter$count = 70171;
	#10 counter$count = 70172;
	#10 counter$count = 70173;
	#10 counter$count = 70174;
	#10 counter$count = 70175;
	#10 counter$count = 70176;
	#10 counter$count = 70177;
	#10 counter$count = 70178;
	#10 counter$count = 70179;
	#10 counter$count = 70180;
	#10 counter$count = 70181;
	#10 counter$count = 70182;
	#10 counter$count = 70183;
	#10 counter$count = 70184;
	#10 counter$count = 70185;
	#10 counter$count = 70186;
	#10 counter$count = 70187;
	#10 counter$count = 70188;
	#10 counter$count = 70189;
	#10 counter$count = 70190;
	#10 counter$count = 70191;
	#10 counter$count = 70192;
	#10 counter$count = 70193;
	#10 counter$count = 70194;
	#10 counter$count = 70195;
	#10 counter$count = 70196;
	#10 counter$count = 70197;
	#10 counter$count = 70198;
	#10 counter$count = 70199;
	#10 counter$count = 70200;
	#10 counter$count = 70201;
	#10 counter$count = 70202;
	#10 counter$count = 70203;
	#10 counter$count = 70204;
	#10 counter$count = 70205;
	#10 counter$count = 70206;
	#10 counter$count = 70207;
	#10 counter$count = 70208;
	#10 counter$count = 70209;
	#10 counter$count = 70210;
	#10 counter$count = 70211;
	#10 counter$count = 70212;
	#10 counter$count = 70213;
	#10 counter$count = 70214;
	#10 counter$count = 70215;
	#10 counter$count = 70216;
	#10 counter$count = 70217;
	#10 counter$count = 70218;
	#10 counter$count = 70219;
	#10 counter$count = 70220;
	#10 counter$count = 70221;
	#10 counter$count = 70222;
	#10 counter$count = 70223;
	#10 counter$count = 70224;
	#10 counter$count = 70225;
	#10 counter$count = 70226;
	#10 counter$count = 70227;
	#10 counter$count = 70228;
	#10 counter$count = 70229;
	#10 counter$count = 70230;
	#10 counter$count = 70231;
	#10 counter$count = 70232;
	#10 counter$count = 70233;
	#10 counter$count = 70234;
	#10 counter$count = 70235;
	#10 counter$count = 70236;
	#10 counter$count = 70237;
	#10 counter$count = 70238;
	#10 counter$count = 70239;
	#10 counter$count = 70240;
	#10 counter$count = 70241;
	#10 counter$count = 70242;
	#10 counter$count = 70243;
	#10 counter$count = 70244;
	#10 counter$count = 70245;
	#10 counter$count = 70246;
	#10 counter$count = 70247;
	#10 counter$count = 70248;
	#10 counter$count = 70249;
	#10 counter$count = 70250;
	#10 counter$count = 70251;
	#10 counter$count = 70252;
	#10 counter$count = 70253;
	#10 counter$count = 70254;
	#10 counter$count = 70255;
	#10 counter$count = 70256;
	#10 counter$count = 70257;
	#10 counter$count = 70258;
	#10 counter$count = 70259;
	#10 counter$count = 70260;
	#10 counter$count = 70261;
	#10 counter$count = 70262;
	#10 counter$count = 70263;
	#10 counter$count = 70264;
	#10 counter$count = 70265;
	#10 counter$count = 70266;
	#10 counter$count = 70267;
	#10 counter$count = 70268;
	#10 counter$count = 70269;
	#10 counter$count = 70270;
	#10 counter$count = 70271;
	#10 counter$count = 70272;
	#10 counter$count = 70273;
	#10 counter$count = 70274;
	#10 counter$count = 70275;
	#10 counter$count = 70276;
	#10 counter$count = 70277;
	#10 counter$count = 70278;
	#10 counter$count = 70279;
	#10 counter$count = 70280;
	#10 counter$count = 70281;
	#10 counter$count = 70282;
	#10 counter$count = 70283;
	#10 counter$count = 70284;
	#10 counter$count = 70285;
	#10 counter$count = 70286;
	#10 counter$count = 70287;
	#10 counter$count = 70288;
	#10 counter$count = 70289;
	#10 counter$count = 70290;
	#10 counter$count = 70291;
	#10 counter$count = 70292;
	#10 counter$count = 70293;
	#10 counter$count = 70294;
	#10 counter$count = 70295;
	#10 counter$count = 70296;
	#10 counter$count = 70297;
	#10 counter$count = 70298;
	#10 counter$count = 70299;
	#10 counter$count = 70300;
	#10 counter$count = 70301;
	#10 counter$count = 70302;
	#10 counter$count = 70303;
	#10 counter$count = 70304;
	#10 counter$count = 70305;
	#10 counter$count = 70306;
	#10 counter$count = 70307;
	#10 counter$count = 70308;
	#10 counter$count = 70309;
	#10 counter$count = 70310;
	#10 counter$count = 70311;
	#10 counter$count = 70312;
	#10 counter$count = 70313;
	#10 counter$count = 70314;
	#10 counter$count = 70315;
	#10 counter$count = 70316;
	#10 counter$count = 70317;
	#10 counter$count = 70318;
	#10 counter$count = 70319;
	#10 counter$count = 70320;
	#10 counter$count = 70321;
	#10 counter$count = 70322;
	#10 counter$count = 70323;
	#10 counter$count = 70324;
	#10 counter$count = 70325;
	#10 counter$count = 70326;
	#10 counter$count = 70327;
	#10 counter$count = 70328;
	#10 counter$count = 70329;
	#10 counter$count = 70330;
	#10 counter$count = 70331;
	#10 counter$count = 70332;
	#10 counter$count = 70333;
	#10 counter$count = 70334;
	#10 counter$count = 70335;
	#10 counter$count = 70336;
	#10 counter$count = 70337;
	#10 counter$count = 70338;
	#10 counter$count = 70339;
	#10 counter$count = 70340;
	#10 counter$count = 70341;
	#10 counter$count = 70342;
	#10 counter$count = 70343;
	#10 counter$count = 70344;
	#10 counter$count = 70345;
	#10 counter$count = 70346;
	#10 counter$count = 70347;
	#10 counter$count = 70348;
	#10 counter$count = 70349;
	#10 counter$count = 70350;
	#10 counter$count = 70351;
	#10 counter$count = 70352;
	#10 counter$count = 70353;
	#10 counter$count = 70354;
	#10 counter$count = 70355;
	#10 counter$count = 70356;
	#10 counter$count = 70357;
	#10 counter$count = 70358;
	#10 counter$count = 70359;
	#10 counter$count = 70360;
	#10 counter$count = 70361;
	#10 counter$count = 70362;
	#10 counter$count = 70363;
	#10 counter$count = 70364;
	#10 counter$count = 70365;
	#10 counter$count = 70366;
	#10 counter$count = 70367;
	#10 counter$count = 70368;
	#10 counter$count = 70369;
	#10 counter$count = 70370;
	#10 counter$count = 70371;
	#10 counter$count = 70372;
	#10 counter$count = 70373;
	#10 counter$count = 70374;
	#10 counter$count = 70375;
	#10 counter$count = 70376;
	#10 counter$count = 70377;
	#10 counter$count = 70378;
	#10 counter$count = 70379;
	#10 counter$count = 70380;
	#10 counter$count = 70381;
	#10 counter$count = 70382;
	#10 counter$count = 70383;
	#10 counter$count = 70384;
	#10 counter$count = 70385;
	#10 counter$count = 70386;
	#10 counter$count = 70387;
	#10 counter$count = 70388;
	#10 counter$count = 70389;
	#10 counter$count = 70390;
	#10 counter$count = 70391;
	#10 counter$count = 70392;
	#10 counter$count = 70393;
	#10 counter$count = 70394;
	#10 counter$count = 70395;
	#10 counter$count = 70396;
	#10 counter$count = 70397;
	#10 counter$count = 70398;
	#10 counter$count = 70399;
	#10 counter$count = 70400;
	#10 counter$count = 70401;
	#10 counter$count = 70402;
	#10 counter$count = 70403;
	#10 counter$count = 70404;
	#10 counter$count = 70405;
	#10 counter$count = 70406;
	#10 counter$count = 70407;
	#10 counter$count = 70408;
	#10 counter$count = 70409;
	#10 counter$count = 70410;
	#10 counter$count = 70411;
	#10 counter$count = 70412;
	#10 counter$count = 70413;
	#10 counter$count = 70414;
	#10 counter$count = 70415;
	#10 counter$count = 70416;
	#10 counter$count = 70417;
	#10 counter$count = 70418;
	#10 counter$count = 70419;
	#10 counter$count = 70420;
	#10 counter$count = 70421;
	#10 counter$count = 70422;
	#10 counter$count = 70423;
	#10 counter$count = 70424;
	#10 counter$count = 70425;
	#10 counter$count = 70426;
	#10 counter$count = 70427;
	#10 counter$count = 70428;
	#10 counter$count = 70429;
	#10 counter$count = 70430;
	#10 counter$count = 70431;
	#10 counter$count = 70432;
	#10 counter$count = 70433;
	#10 counter$count = 70434;
	#10 counter$count = 70435;
	#10 counter$count = 70436;
	#10 counter$count = 70437;
	#10 counter$count = 70438;
	#10 counter$count = 70439;
	#10 counter$count = 70440;
	#10 counter$count = 70441;
	#10 counter$count = 70442;
	#10 counter$count = 70443;
	#10 counter$count = 70444;
	#10 counter$count = 70445;
	#10 counter$count = 70446;
	#10 counter$count = 70447;
	#10 counter$count = 70448;
	#10 counter$count = 70449;
	#10 counter$count = 70450;
	#10 counter$count = 70451;
	#10 counter$count = 70452;
	#10 counter$count = 70453;
	#10 counter$count = 70454;
	#10 counter$count = 70455;
	#10 counter$count = 70456;
	#10 counter$count = 70457;
	#10 counter$count = 70458;
	#10 counter$count = 70459;
	#10 counter$count = 70460;
	#10 counter$count = 70461;
	#10 counter$count = 70462;
	#10 counter$count = 70463;
	#10 counter$count = 70464;
	#10 counter$count = 70465;
	#10 counter$count = 70466;
	#10 counter$count = 70467;
	#10 counter$count = 70468;
	#10 counter$count = 70469;
	#10 counter$count = 70470;
	#10 counter$count = 70471;
	#10 counter$count = 70472;
	#10 counter$count = 70473;
	#10 counter$count = 70474;
	#10 counter$count = 70475;
	#10 counter$count = 70476;
	#10 counter$count = 70477;
	#10 counter$count = 70478;
	#10 counter$count = 70479;
	#10 counter$count = 70480;
	#10 counter$count = 70481;
	#10 counter$count = 70482;
	#10 counter$count = 70483;
	#10 counter$count = 70484;
	#10 counter$count = 70485;
	#10 counter$count = 70486;
	#10 counter$count = 70487;
	#10 counter$count = 70488;
	#10 counter$count = 70489;
	#10 counter$count = 70490;
	#10 counter$count = 70491;
	#10 counter$count = 70492;
	#10 counter$count = 70493;
	#10 counter$count = 70494;
	#10 counter$count = 70495;
	#10 counter$count = 70496;
	#10 counter$count = 70497;
	#10 counter$count = 70498;
	#10 counter$count = 70499;
	#10 counter$count = 70500;
	#10 counter$count = 70501;
	#10 counter$count = 70502;
	#10 counter$count = 70503;
	#10 counter$count = 70504;
	#10 counter$count = 70505;
	#10 counter$count = 70506;
	#10 counter$count = 70507;
	#10 counter$count = 70508;
	#10 counter$count = 70509;
	#10 counter$count = 70510;
	#10 counter$count = 70511;
	#10 counter$count = 70512;
	#10 counter$count = 70513;
	#10 counter$count = 70514;
	#10 counter$count = 70515;
	#10 counter$count = 70516;
	#10 counter$count = 70517;
	#10 counter$count = 70518;
	#10 counter$count = 70519;
	#10 counter$count = 70520;
	#10 counter$count = 70521;
	#10 counter$count = 70522;
	#10 counter$count = 70523;
	#10 counter$count = 70524;
	#10 counter$count = 70525;
	#10 counter$count = 70526;
	#10 counter$count = 70527;
	#10 counter$count = 70528;
	#10 counter$count = 70529;
	#10 counter$count = 70530;
	#10 counter$count = 70531;
	#10 counter$count = 70532;
	#10 counter$count = 70533;
	#10 counter$count = 70534;
	#10 counter$count = 70535;
	#10 counter$count = 70536;
	#10 counter$count = 70537;
	#10 counter$count = 70538;
	#10 counter$count = 70539;
	#10 counter$count = 70540;
	#10 counter$count = 70541;
	#10 counter$count = 70542;
	#10 counter$count = 70543;
	#10 counter$count = 70544;
	#10 counter$count = 70545;
	#10 counter$count = 70546;
	#10 counter$count = 70547;
	#10 counter$count = 70548;
	#10 counter$count = 70549;
	#10 counter$count = 70550;
	#10 counter$count = 70551;
	#10 counter$count = 70552;
	#10 counter$count = 70553;
	#10 counter$count = 70554;
	#10 counter$count = 70555;
	#10 counter$count = 70556;
	#10 counter$count = 70557;
	#10 counter$count = 70558;
	#10 counter$count = 70559;
	#10 counter$count = 70560;
	#10 counter$count = 70561;
	#10 counter$count = 70562;
	#10 counter$count = 70563;
	#10 counter$count = 70564;
	#10 counter$count = 70565;
	#10 counter$count = 70566;
	#10 counter$count = 70567;
	#10 counter$count = 70568;
	#10 counter$count = 70569;
	#10 counter$count = 70570;
	#10 counter$count = 70571;
	#10 counter$count = 70572;
	#10 counter$count = 70573;
	#10 counter$count = 70574;
	#10 counter$count = 70575;
	#10 counter$count = 70576;
	#10 counter$count = 70577;
	#10 counter$count = 70578;
	#10 counter$count = 70579;
	#10 counter$count = 70580;
	#10 counter$count = 70581;
	#10 counter$count = 70582;
	#10 counter$count = 70583;
	#10 counter$count = 70584;
	#10 counter$count = 70585;
	#10 counter$count = 70586;
	#10 counter$count = 70587;
	#10 counter$count = 70588;
	#10 counter$count = 70589;
	#10 counter$count = 70590;
	#10 counter$count = 70591;
	#10 counter$count = 70592;
	#10 counter$count = 70593;
	#10 counter$count = 70594;
	#10 counter$count = 70595;
	#10 counter$count = 70596;
	#10 counter$count = 70597;
	#10 counter$count = 70598;
	#10 counter$count = 70599;
	#10 counter$count = 70600;
	#10 counter$count = 70601;
	#10 counter$count = 70602;
	#10 counter$count = 70603;
	#10 counter$count = 70604;
	#10 counter$count = 70605;
	#10 counter$count = 70606;
	#10 counter$count = 70607;
	#10 counter$count = 70608;
	#10 counter$count = 70609;
	#10 counter$count = 70610;
	#10 counter$count = 70611;
	#10 counter$count = 70612;
	#10 counter$count = 70613;
	#10 counter$count = 70614;
	#10 counter$count = 70615;
	#10 counter$count = 70616;
	#10 counter$count = 70617;
	#10 counter$count = 70618;
	#10 counter$count = 70619;
	#10 counter$count = 70620;
	#10 counter$count = 70621;
	#10 counter$count = 70622;
	#10 counter$count = 70623;
	#10 counter$count = 70624;
	#10 counter$count = 70625;
	#10 counter$count = 70626;
	#10 counter$count = 70627;
	#10 counter$count = 70628;
	#10 counter$count = 70629;
	#10 counter$count = 70630;
	#10 counter$count = 70631;
	#10 counter$count = 70632;
	#10 counter$count = 70633;
	#10 counter$count = 70634;
	#10 counter$count = 70635;
	#10 counter$count = 70636;
	#10 counter$count = 70637;
	#10 counter$count = 70638;
	#10 counter$count = 70639;
	#10 counter$count = 70640;
	#10 counter$count = 70641;
	#10 counter$count = 70642;
	#10 counter$count = 70643;
	#10 counter$count = 70644;
	#10 counter$count = 70645;
	#10 counter$count = 70646;
	#10 counter$count = 70647;
	#10 counter$count = 70648;
	#10 counter$count = 70649;
	#10 counter$count = 70650;
	#10 counter$count = 70651;
	#10 counter$count = 70652;
	#10 counter$count = 70653;
	#10 counter$count = 70654;
	#10 counter$count = 70655;
	#10 counter$count = 70656;
	#10 counter$count = 70657;
	#10 counter$count = 70658;
	#10 counter$count = 70659;
	#10 counter$count = 70660;
	#10 counter$count = 70661;
	#10 counter$count = 70662;
	#10 counter$count = 70663;
	#10 counter$count = 70664;
	#10 counter$count = 70665;
	#10 counter$count = 70666;
	#10 counter$count = 70667;
	#10 counter$count = 70668;
	#10 counter$count = 70669;
	#10 counter$count = 70670;
	#10 counter$count = 70671;
	#10 counter$count = 70672;
	#10 counter$count = 70673;
	#10 counter$count = 70674;
	#10 counter$count = 70675;
	#10 counter$count = 70676;
	#10 counter$count = 70677;
	#10 counter$count = 70678;
	#10 counter$count = 70679;
	#10 counter$count = 70680;
	#10 counter$count = 70681;
	#10 counter$count = 70682;
	#10 counter$count = 70683;
	#10 counter$count = 70684;
	#10 counter$count = 70685;
	#10 counter$count = 70686;
	#10 counter$count = 70687;
	#10 counter$count = 70688;
	#10 counter$count = 70689;
	#10 counter$count = 70690;
	#10 counter$count = 70691;
	#10 counter$count = 70692;
	#10 counter$count = 70693;
	#10 counter$count = 70694;
	#10 counter$count = 70695;
	#10 counter$count = 70696;
	#10 counter$count = 70697;
	#10 counter$count = 70698;
	#10 counter$count = 70699;
	#10 counter$count = 70700;
	#10 counter$count = 70701;
	#10 counter$count = 70702;
	#10 counter$count = 70703;
	#10 counter$count = 70704;
	#10 counter$count = 70705;
	#10 counter$count = 70706;
	#10 counter$count = 70707;
	#10 counter$count = 70708;
	#10 counter$count = 70709;
	#10 counter$count = 70710;
	#10 counter$count = 70711;
	#10 counter$count = 70712;
	#10 counter$count = 70713;
	#10 counter$count = 70714;
	#10 counter$count = 70715;
	#10 counter$count = 70716;
	#10 counter$count = 70717;
	#10 counter$count = 70718;
	#10 counter$count = 70719;
	#10 counter$count = 70720;
	#10 counter$count = 70721;
	#10 counter$count = 70722;
	#10 counter$count = 70723;
	#10 counter$count = 70724;
	#10 counter$count = 70725;
	#10 counter$count = 70726;
	#10 counter$count = 70727;
	#10 counter$count = 70728;
	#10 counter$count = 70729;
	#10 counter$count = 70730;
	#10 counter$count = 70731;
	#10 counter$count = 70732;
	#10 counter$count = 70733;
	#10 counter$count = 70734;
	#10 counter$count = 70735;
	#10 counter$count = 70736;
	#10 counter$count = 70737;
	#10 counter$count = 70738;
	#10 counter$count = 70739;
	#10 counter$count = 70740;
	#10 counter$count = 70741;
	#10 counter$count = 70742;
	#10 counter$count = 70743;
	#10 counter$count = 70744;
	#10 counter$count = 70745;
	#10 counter$count = 70746;
	#10 counter$count = 70747;
	#10 counter$count = 70748;
	#10 counter$count = 70749;
	#10 counter$count = 70750;
	#10 counter$count = 70751;
	#10 counter$count = 70752;
	#10 counter$count = 70753;
	#10 counter$count = 70754;
	#10 counter$count = 70755;
	#10 counter$count = 70756;
	#10 counter$count = 70757;
	#10 counter$count = 70758;
	#10 counter$count = 70759;
	#10 counter$count = 70760;
	#10 counter$count = 70761;
	#10 counter$count = 70762;
	#10 counter$count = 70763;
	#10 counter$count = 70764;
	#10 counter$count = 70765;
	#10 counter$count = 70766;
	#10 counter$count = 70767;
	#10 counter$count = 70768;
	#10 counter$count = 70769;
	#10 counter$count = 70770;
	#10 counter$count = 70771;
	#10 counter$count = 70772;
	#10 counter$count = 70773;
	#10 counter$count = 70774;
	#10 counter$count = 70775;
	#10 counter$count = 70776;
	#10 counter$count = 70777;
	#10 counter$count = 70778;
	#10 counter$count = 70779;
	#10 counter$count = 70780;
	#10 counter$count = 70781;
	#10 counter$count = 70782;
	#10 counter$count = 70783;
	#10 counter$count = 70784;
	#10 counter$count = 70785;
	#10 counter$count = 70786;
	#10 counter$count = 70787;
	#10 counter$count = 70788;
	#10 counter$count = 70789;
	#10 counter$count = 70790;
	#10 counter$count = 70791;
	#10 counter$count = 70792;
	#10 counter$count = 70793;
	#10 counter$count = 70794;
	#10 counter$count = 70795;
	#10 counter$count = 70796;
	#10 counter$count = 70797;
	#10 counter$count = 70798;
	#10 counter$count = 70799;
	#10 counter$count = 70800;
	#10 counter$count = 70801;
	#10 counter$count = 70802;
	#10 counter$count = 70803;
	#10 counter$count = 70804;
	#10 counter$count = 70805;
	#10 counter$count = 70806;
	#10 counter$count = 70807;
	#10 counter$count = 70808;
	#10 counter$count = 70809;
	#10 counter$count = 70810;
	#10 counter$count = 70811;
	#10 counter$count = 70812;
	#10 counter$count = 70813;
	#10 counter$count = 70814;
	#10 counter$count = 70815;
	#10 counter$count = 70816;
	#10 counter$count = 70817;
	#10 counter$count = 70818;
	#10 counter$count = 70819;
	#10 counter$count = 70820;
	#10 counter$count = 70821;
	#10 counter$count = 70822;
	#10 counter$count = 70823;
	#10 counter$count = 70824;
	#10 counter$count = 70825;
	#10 counter$count = 70826;
	#10 counter$count = 70827;
	#10 counter$count = 70828;
	#10 counter$count = 70829;
	#10 counter$count = 70830;
	#10 counter$count = 70831;
	#10 counter$count = 70832;
	#10 counter$count = 70833;
	#10 counter$count = 70834;
	#10 counter$count = 70835;
	#10 counter$count = 70836;
	#10 counter$count = 70837;
	#10 counter$count = 70838;
	#10 counter$count = 70839;
	#10 counter$count = 70840;
	#10 counter$count = 70841;
	#10 counter$count = 70842;
	#10 counter$count = 70843;
	#10 counter$count = 70844;
	#10 counter$count = 70845;
	#10 counter$count = 70846;
	#10 counter$count = 70847;
	#10 counter$count = 70848;
	#10 counter$count = 70849;
	#10 counter$count = 70850;
	#10 counter$count = 70851;
	#10 counter$count = 70852;
	#10 counter$count = 70853;
	#10 counter$count = 70854;
	#10 counter$count = 70855;
	#10 counter$count = 70856;
	#10 counter$count = 70857;
	#10 counter$count = 70858;
	#10 counter$count = 70859;
	#10 counter$count = 70860;
	#10 counter$count = 70861;
	#10 counter$count = 70862;
	#10 counter$count = 70863;
	#10 counter$count = 70864;
	#10 counter$count = 70865;
	#10 counter$count = 70866;
	#10 counter$count = 70867;
	#10 counter$count = 70868;
	#10 counter$count = 70869;
	#10 counter$count = 70870;
	#10 counter$count = 70871;
	#10 counter$count = 70872;
	#10 counter$count = 70873;
	#10 counter$count = 70874;
	#10 counter$count = 70875;
	#10 counter$count = 70876;
	#10 counter$count = 70877;
	#10 counter$count = 70878;
	#10 counter$count = 70879;
	#10 counter$count = 70880;
	#10 counter$count = 70881;
	#10 counter$count = 70882;
	#10 counter$count = 70883;
	#10 counter$count = 70884;
	#10 counter$count = 70885;
	#10 counter$count = 70886;
	#10 counter$count = 70887;
	#10 counter$count = 70888;
	#10 counter$count = 70889;
	#10 counter$count = 70890;
	#10 counter$count = 70891;
	#10 counter$count = 70892;
	#10 counter$count = 70893;
	#10 counter$count = 70894;
	#10 counter$count = 70895;
	#10 counter$count = 70896;
	#10 counter$count = 70897;
	#10 counter$count = 70898;
	#10 counter$count = 70899;
	#10 counter$count = 70900;
	#10 counter$count = 70901;
	#10 counter$count = 70902;
	#10 counter$count = 70903;
	#10 counter$count = 70904;
	#10 counter$count = 70905;
	#10 counter$count = 70906;
	#10 counter$count = 70907;
	#10 counter$count = 70908;
	#10 counter$count = 70909;
	#10 counter$count = 70910;
	#10 counter$count = 70911;
	#10 counter$count = 70912;
	#10 counter$count = 70913;
	#10 counter$count = 70914;
	#10 counter$count = 70915;
	#10 counter$count = 70916;
	#10 counter$count = 70917;
	#10 counter$count = 70918;
	#10 counter$count = 70919;
	#10 counter$count = 70920;
	#10 counter$count = 70921;
	#10 counter$count = 70922;
	#10 counter$count = 70923;
	#10 counter$count = 70924;
	#10 counter$count = 70925;
	#10 counter$count = 70926;
	#10 counter$count = 70927;
	#10 counter$count = 70928;
	#10 counter$count = 70929;
	#10 counter$count = 70930;
	#10 counter$count = 70931;
	#10 counter$count = 70932;
	#10 counter$count = 70933;
	#10 counter$count = 70934;
	#10 counter$count = 70935;
	#10 counter$count = 70936;
	#10 counter$count = 70937;
	#10 counter$count = 70938;
	#10 counter$count = 70939;
	#10 counter$count = 70940;
	#10 counter$count = 70941;
	#10 counter$count = 70942;
	#10 counter$count = 70943;
	#10 counter$count = 70944;
	#10 counter$count = 70945;
	#10 counter$count = 70946;
	#10 counter$count = 70947;
	#10 counter$count = 70948;
	#10 counter$count = 70949;
	#10 counter$count = 70950;
	#10 counter$count = 70951;
	#10 counter$count = 70952;
	#10 counter$count = 70953;
	#10 counter$count = 70954;
	#10 counter$count = 70955;
	#10 counter$count = 70956;
	#10 counter$count = 70957;
	#10 counter$count = 70958;
	#10 counter$count = 70959;
	#10 counter$count = 70960;
	#10 counter$count = 70961;
	#10 counter$count = 70962;
	#10 counter$count = 70963;
	#10 counter$count = 70964;
	#10 counter$count = 70965;
	#10 counter$count = 70966;
	#10 counter$count = 70967;
	#10 counter$count = 70968;
	#10 counter$count = 70969;
	#10 counter$count = 70970;
	#10 counter$count = 70971;
	#10 counter$count = 70972;
	#10 counter$count = 70973;
	#10 counter$count = 70974;
	#10 counter$count = 70975;
	#10 counter$count = 70976;
	#10 counter$count = 70977;
	#10 counter$count = 70978;
	#10 counter$count = 70979;
	#10 counter$count = 70980;
	#10 counter$count = 70981;
	#10 counter$count = 70982;
	#10 counter$count = 70983;
	#10 counter$count = 70984;
	#10 counter$count = 70985;
	#10 counter$count = 70986;
	#10 counter$count = 70987;
	#10 counter$count = 70988;
	#10 counter$count = 70989;
	#10 counter$count = 70990;
	#10 counter$count = 70991;
	#10 counter$count = 70992;
	#10 counter$count = 70993;
	#10 counter$count = 70994;
	#10 counter$count = 70995;
	#10 counter$count = 70996;
	#10 counter$count = 70997;
	#10 counter$count = 70998;
	#10 counter$count = 70999;
	#10 counter$count = 71000;
	#10 counter$count = 71001;
	#10 counter$count = 71002;
	#10 counter$count = 71003;
	#10 counter$count = 71004;
	#10 counter$count = 71005;
	#10 counter$count = 71006;
	#10 counter$count = 71007;
	#10 counter$count = 71008;
	#10 counter$count = 71009;
	#10 counter$count = 71010;
	#10 counter$count = 71011;
	#10 counter$count = 71012;
	#10 counter$count = 71013;
	#10 counter$count = 71014;
	#10 counter$count = 71015;
	#10 counter$count = 71016;
	#10 counter$count = 71017;
	#10 counter$count = 71018;
	#10 counter$count = 71019;
	#10 counter$count = 71020;
	#10 counter$count = 71021;
	#10 counter$count = 71022;
	#10 counter$count = 71023;
	#10 counter$count = 71024;
	#10 counter$count = 71025;
	#10 counter$count = 71026;
	#10 counter$count = 71027;
	#10 counter$count = 71028;
	#10 counter$count = 71029;
	#10 counter$count = 71030;
	#10 counter$count = 71031;
	#10 counter$count = 71032;
	#10 counter$count = 71033;
	#10 counter$count = 71034;
	#10 counter$count = 71035;
	#10 counter$count = 71036;
	#10 counter$count = 71037;
	#10 counter$count = 71038;
	#10 counter$count = 71039;
	#10 counter$count = 71040;
	#10 counter$count = 71041;
	#10 counter$count = 71042;
	#10 counter$count = 71043;
	#10 counter$count = 71044;
	#10 counter$count = 71045;
	#10 counter$count = 71046;
	#10 counter$count = 71047;
	#10 counter$count = 71048;
	#10 counter$count = 71049;
	#10 counter$count = 71050;
	#10 counter$count = 71051;
	#10 counter$count = 71052;
	#10 counter$count = 71053;
	#10 counter$count = 71054;
	#10 counter$count = 71055;
	#10 counter$count = 71056;
	#10 counter$count = 71057;
	#10 counter$count = 71058;
	#10 counter$count = 71059;
	#10 counter$count = 71060;
	#10 counter$count = 71061;
	#10 counter$count = 71062;
	#10 counter$count = 71063;
	#10 counter$count = 71064;
	#10 counter$count = 71065;
	#10 counter$count = 71066;
	#10 counter$count = 71067;
	#10 counter$count = 71068;
	#10 counter$count = 71069;
	#10 counter$count = 71070;
	#10 counter$count = 71071;
	#10 counter$count = 71072;
	#10 counter$count = 71073;
	#10 counter$count = 71074;
	#10 counter$count = 71075;
	#10 counter$count = 71076;
	#10 counter$count = 71077;
	#10 counter$count = 71078;
	#10 counter$count = 71079;
	#10 counter$count = 71080;
	#10 counter$count = 71081;
	#10 counter$count = 71082;
	#10 counter$count = 71083;
	#10 counter$count = 71084;
	#10 counter$count = 71085;
	#10 counter$count = 71086;
	#10 counter$count = 71087;
	#10 counter$count = 71088;
	#10 counter$count = 71089;
	#10 counter$count = 71090;
	#10 counter$count = 71091;
	#10 counter$count = 71092;
	#10 counter$count = 71093;
	#10 counter$count = 71094;
	#10 counter$count = 71095;
	#10 counter$count = 71096;
	#10 counter$count = 71097;
	#10 counter$count = 71098;
	#10 counter$count = 71099;
	#10 counter$count = 71100;
	#10 counter$count = 71101;
	#10 counter$count = 71102;
	#10 counter$count = 71103;
	#10 counter$count = 71104;
	#10 counter$count = 71105;
	#10 counter$count = 71106;
	#10 counter$count = 71107;
	#10 counter$count = 71108;
	#10 counter$count = 71109;
	#10 counter$count = 71110;
	#10 counter$count = 71111;
	#10 counter$count = 71112;
	#10 counter$count = 71113;
	#10 counter$count = 71114;
	#10 counter$count = 71115;
	#10 counter$count = 71116;
	#10 counter$count = 71117;
	#10 counter$count = 71118;
	#10 counter$count = 71119;
	#10 counter$count = 71120;
	#10 counter$count = 71121;
	#10 counter$count = 71122;
	#10 counter$count = 71123;
	#10 counter$count = 71124;
	#10 counter$count = 71125;
	#10 counter$count = 71126;
	#10 counter$count = 71127;
	#10 counter$count = 71128;
	#10 counter$count = 71129;
	#10 counter$count = 71130;
	#10 counter$count = 71131;
	#10 counter$count = 71132;
	#10 counter$count = 71133;
	#10 counter$count = 71134;
	#10 counter$count = 71135;
	#10 counter$count = 71136;
	#10 counter$count = 71137;
	#10 counter$count = 71138;
	#10 counter$count = 71139;
	#10 counter$count = 71140;
	#10 counter$count = 71141;
	#10 counter$count = 71142;
	#10 counter$count = 71143;
	#10 counter$count = 71144;
	#10 counter$count = 71145;
	#10 counter$count = 71146;
	#10 counter$count = 71147;
	#10 counter$count = 71148;
	#10 counter$count = 71149;
	#10 counter$count = 71150;
	#10 counter$count = 71151;
	#10 counter$count = 71152;
	#10 counter$count = 71153;
	#10 counter$count = 71154;
	#10 counter$count = 71155;
	#10 counter$count = 71156;
	#10 counter$count = 71157;
	#10 counter$count = 71158;
	#10 counter$count = 71159;
	#10 counter$count = 71160;
	#10 counter$count = 71161;
	#10 counter$count = 71162;
	#10 counter$count = 71163;
	#10 counter$count = 71164;
	#10 counter$count = 71165;
	#10 counter$count = 71166;
	#10 counter$count = 71167;
	#10 counter$count = 71168;
	#10 counter$count = 71169;
	#10 counter$count = 71170;
	#10 counter$count = 71171;
	#10 counter$count = 71172;
	#10 counter$count = 71173;
	#10 counter$count = 71174;
	#10 counter$count = 71175;
	#10 counter$count = 71176;
	#10 counter$count = 71177;
	#10 counter$count = 71178;
	#10 counter$count = 71179;
	#10 counter$count = 71180;
	#10 counter$count = 71181;
	#10 counter$count = 71182;
	#10 counter$count = 71183;
	#10 counter$count = 71184;
	#10 counter$count = 71185;
	#10 counter$count = 71186;
	#10 counter$count = 71187;
	#10 counter$count = 71188;
	#10 counter$count = 71189;
	#10 counter$count = 71190;
	#10 counter$count = 71191;
	#10 counter$count = 71192;
	#10 counter$count = 71193;
	#10 counter$count = 71194;
	#10 counter$count = 71195;
	#10 counter$count = 71196;
	#10 counter$count = 71197;
	#10 counter$count = 71198;
	#10 counter$count = 71199;
	#10 counter$count = 71200;
	#10 counter$count = 71201;
	#10 counter$count = 71202;
	#10 counter$count = 71203;
	#10 counter$count = 71204;
	#10 counter$count = 71205;
	#10 counter$count = 71206;
	#10 counter$count = 71207;
	#10 counter$count = 71208;
	#10 counter$count = 71209;
	#10 counter$count = 71210;
	#10 counter$count = 71211;
	#10 counter$count = 71212;
	#10 counter$count = 71213;
	#10 counter$count = 71214;
	#10 counter$count = 71215;
	#10 counter$count = 71216;
	#10 counter$count = 71217;
	#10 counter$count = 71218;
	#10 counter$count = 71219;
	#10 counter$count = 71220;
	#10 counter$count = 71221;
	#10 counter$count = 71222;
	#10 counter$count = 71223;
	#10 counter$count = 71224;
	#10 counter$count = 71225;
	#10 counter$count = 71226;
	#10 counter$count = 71227;
	#10 counter$count = 71228;
	#10 counter$count = 71229;
	#10 counter$count = 71230;
	#10 counter$count = 71231;
	#10 counter$count = 71232;
	#10 counter$count = 71233;
	#10 counter$count = 71234;
	#10 counter$count = 71235;
	#10 counter$count = 71236;
	#10 counter$count = 71237;
	#10 counter$count = 71238;
	#10 counter$count = 71239;
	#10 counter$count = 71240;
	#10 counter$count = 71241;
	#10 counter$count = 71242;
	#10 counter$count = 71243;
	#10 counter$count = 71244;
	#10 counter$count = 71245;
	#10 counter$count = 71246;
	#10 counter$count = 71247;
	#10 counter$count = 71248;
	#10 counter$count = 71249;
	#10 counter$count = 71250;
	#10 counter$count = 71251;
	#10 counter$count = 71252;
	#10 counter$count = 71253;
	#10 counter$count = 71254;
	#10 counter$count = 71255;
	#10 counter$count = 71256;
	#10 counter$count = 71257;
	#10 counter$count = 71258;
	#10 counter$count = 71259;
	#10 counter$count = 71260;
	#10 counter$count = 71261;
	#10 counter$count = 71262;
	#10 counter$count = 71263;
	#10 counter$count = 71264;
	#10 counter$count = 71265;
	#10 counter$count = 71266;
	#10 counter$count = 71267;
	#10 counter$count = 71268;
	#10 counter$count = 71269;
	#10 counter$count = 71270;
	#10 counter$count = 71271;
	#10 counter$count = 71272;
	#10 counter$count = 71273;
	#10 counter$count = 71274;
	#10 counter$count = 71275;
	#10 counter$count = 71276;
	#10 counter$count = 71277;
	#10 counter$count = 71278;
	#10 counter$count = 71279;
	#10 counter$count = 71280;
	#10 counter$count = 71281;
	#10 counter$count = 71282;
	#10 counter$count = 71283;
	#10 counter$count = 71284;
	#10 counter$count = 71285;
	#10 counter$count = 71286;
	#10 counter$count = 71287;
	#10 counter$count = 71288;
	#10 counter$count = 71289;
	#10 counter$count = 71290;
	#10 counter$count = 71291;
	#10 counter$count = 71292;
	#10 counter$count = 71293;
	#10 counter$count = 71294;
	#10 counter$count = 71295;
	#10 counter$count = 71296;
	#10 counter$count = 71297;
	#10 counter$count = 71298;
	#10 counter$count = 71299;
	#10 counter$count = 71300;
	#10 counter$count = 71301;
	#10 counter$count = 71302;
	#10 counter$count = 71303;
	#10 counter$count = 71304;
	#10 counter$count = 71305;
	#10 counter$count = 71306;
	#10 counter$count = 71307;
	#10 counter$count = 71308;
	#10 counter$count = 71309;
	#10 counter$count = 71310;
	#10 counter$count = 71311;
	#10 counter$count = 71312;
	#10 counter$count = 71313;
	#10 counter$count = 71314;
	#10 counter$count = 71315;
	#10 counter$count = 71316;
	#10 counter$count = 71317;
	#10 counter$count = 71318;
	#10 counter$count = 71319;
	#10 counter$count = 71320;
	#10 counter$count = 71321;
	#10 counter$count = 71322;
	#10 counter$count = 71323;
	#10 counter$count = 71324;
	#10 counter$count = 71325;
	#10 counter$count = 71326;
	#10 counter$count = 71327;
	#10 counter$count = 71328;
	#10 counter$count = 71329;
	#10 counter$count = 71330;
	#10 counter$count = 71331;
	#10 counter$count = 71332;
	#10 counter$count = 71333;
	#10 counter$count = 71334;
	#10 counter$count = 71335;
	#10 counter$count = 71336;
	#10 counter$count = 71337;
	#10 counter$count = 71338;
	#10 counter$count = 71339;
	#10 counter$count = 71340;
	#10 counter$count = 71341;
	#10 counter$count = 71342;
	#10 counter$count = 71343;
	#10 counter$count = 71344;
	#10 counter$count = 71345;
	#10 counter$count = 71346;
	#10 counter$count = 71347;
	#10 counter$count = 71348;
	#10 counter$count = 71349;
	#10 counter$count = 71350;
	#10 counter$count = 71351;
	#10 counter$count = 71352;
	#10 counter$count = 71353;
	#10 counter$count = 71354;
	#10 counter$count = 71355;
	#10 counter$count = 71356;
	#10 counter$count = 71357;
	#10 counter$count = 71358;
	#10 counter$count = 71359;
	#10 counter$count = 71360;
	#10 counter$count = 71361;
	#10 counter$count = 71362;
	#10 counter$count = 71363;
	#10 counter$count = 71364;
	#10 counter$count = 71365;
	#10 counter$count = 71366;
	#10 counter$count = 71367;
	#10 counter$count = 71368;
	#10 counter$count = 71369;
	#10 counter$count = 71370;
	#10 counter$count = 71371;
	#10 counter$count = 71372;
	#10 counter$count = 71373;
	#10 counter$count = 71374;
	#10 counter$count = 71375;
	#10 counter$count = 71376;
	#10 counter$count = 71377;
	#10 counter$count = 71378;
	#10 counter$count = 71379;
	#10 counter$count = 71380;
	#10 counter$count = 71381;
	#10 counter$count = 71382;
	#10 counter$count = 71383;
	#10 counter$count = 71384;
	#10 counter$count = 71385;
	#10 counter$count = 71386;
	#10 counter$count = 71387;
	#10 counter$count = 71388;
	#10 counter$count = 71389;
	#10 counter$count = 71390;
	#10 counter$count = 71391;
	#10 counter$count = 71392;
	#10 counter$count = 71393;
	#10 counter$count = 71394;
	#10 counter$count = 71395;
	#10 counter$count = 71396;
	#10 counter$count = 71397;
	#10 counter$count = 71398;
	#10 counter$count = 71399;
	#10 counter$count = 71400;
	#10 counter$count = 71401;
	#10 counter$count = 71402;
	#10 counter$count = 71403;
	#10 counter$count = 71404;
	#10 counter$count = 71405;
	#10 counter$count = 71406;
	#10 counter$count = 71407;
	#10 counter$count = 71408;
	#10 counter$count = 71409;
	#10 counter$count = 71410;
	#10 counter$count = 71411;
	#10 counter$count = 71412;
	#10 counter$count = 71413;
	#10 counter$count = 71414;
	#10 counter$count = 71415;
	#10 counter$count = 71416;
	#10 counter$count = 71417;
	#10 counter$count = 71418;
	#10 counter$count = 71419;
	#10 counter$count = 71420;
	#10 counter$count = 71421;
	#10 counter$count = 71422;
	#10 counter$count = 71423;
	#10 counter$count = 71424;
	#10 counter$count = 71425;
	#10 counter$count = 71426;
	#10 counter$count = 71427;
	#10 counter$count = 71428;
	#10 counter$count = 71429;
	#10 counter$count = 71430;
	#10 counter$count = 71431;
	#10 counter$count = 71432;
	#10 counter$count = 71433;
	#10 counter$count = 71434;
	#10 counter$count = 71435;
	#10 counter$count = 71436;
	#10 counter$count = 71437;
	#10 counter$count = 71438;
	#10 counter$count = 71439;
	#10 counter$count = 71440;
	#10 counter$count = 71441;
	#10 counter$count = 71442;
	#10 counter$count = 71443;
	#10 counter$count = 71444;
	#10 counter$count = 71445;
	#10 counter$count = 71446;
	#10 counter$count = 71447;
	#10 counter$count = 71448;
	#10 counter$count = 71449;
	#10 counter$count = 71450;
	#10 counter$count = 71451;
	#10 counter$count = 71452;
	#10 counter$count = 71453;
	#10 counter$count = 71454;
	#10 counter$count = 71455;
	#10 counter$count = 71456;
	#10 counter$count = 71457;
	#10 counter$count = 71458;
	#10 counter$count = 71459;
	#10 counter$count = 71460;
	#10 counter$count = 71461;
	#10 counter$count = 71462;
	#10 counter$count = 71463;
	#10 counter$count = 71464;
	#10 counter$count = 71465;
	#10 counter$count = 71466;
	#10 counter$count = 71467;
	#10 counter$count = 71468;
	#10 counter$count = 71469;
	#10 counter$count = 71470;
	#10 counter$count = 71471;
	#10 counter$count = 71472;
	#10 counter$count = 71473;
	#10 counter$count = 71474;
	#10 counter$count = 71475;
	#10 counter$count = 71476;
	#10 counter$count = 71477;
	#10 counter$count = 71478;
	#10 counter$count = 71479;
	#10 counter$count = 71480;
	#10 counter$count = 71481;
	#10 counter$count = 71482;
	#10 counter$count = 71483;
	#10 counter$count = 71484;
	#10 counter$count = 71485;
	#10 counter$count = 71486;
	#10 counter$count = 71487;
	#10 counter$count = 71488;
	#10 counter$count = 71489;
	#10 counter$count = 71490;
	#10 counter$count = 71491;
	#10 counter$count = 71492;
	#10 counter$count = 71493;
	#10 counter$count = 71494;
	#10 counter$count = 71495;
	#10 counter$count = 71496;
	#10 counter$count = 71497;
	#10 counter$count = 71498;
	#10 counter$count = 71499;
	#10 counter$count = 71500;
	#10 counter$count = 71501;
	#10 counter$count = 71502;
	#10 counter$count = 71503;
	#10 counter$count = 71504;
	#10 counter$count = 71505;
	#10 counter$count = 71506;
	#10 counter$count = 71507;
	#10 counter$count = 71508;
	#10 counter$count = 71509;
	#10 counter$count = 71510;
	#10 counter$count = 71511;
	#10 counter$count = 71512;
	#10 counter$count = 71513;
	#10 counter$count = 71514;
	#10 counter$count = 71515;
	#10 counter$count = 71516;
	#10 counter$count = 71517;
	#10 counter$count = 71518;
	#10 counter$count = 71519;
	#10 counter$count = 71520;
	#10 counter$count = 71521;
	#10 counter$count = 71522;
	#10 counter$count = 71523;
	#10 counter$count = 71524;
	#10 counter$count = 71525;
	#10 counter$count = 71526;
	#10 counter$count = 71527;
	#10 counter$count = 71528;
	#10 counter$count = 71529;
	#10 counter$count = 71530;
	#10 counter$count = 71531;
	#10 counter$count = 71532;
	#10 counter$count = 71533;
	#10 counter$count = 71534;
	#10 counter$count = 71535;
	#10 counter$count = 71536;
	#10 counter$count = 71537;
	#10 counter$count = 71538;
	#10 counter$count = 71539;
	#10 counter$count = 71540;
	#10 counter$count = 71541;
	#10 counter$count = 71542;
	#10 counter$count = 71543;
	#10 counter$count = 71544;
	#10 counter$count = 71545;
	#10 counter$count = 71546;
	#10 counter$count = 71547;
	#10 counter$count = 71548;
	#10 counter$count = 71549;
	#10 counter$count = 71550;
	#10 counter$count = 71551;
	#10 counter$count = 71552;
	#10 counter$count = 71553;
	#10 counter$count = 71554;
	#10 counter$count = 71555;
	#10 counter$count = 71556;
	#10 counter$count = 71557;
	#10 counter$count = 71558;
	#10 counter$count = 71559;
	#10 counter$count = 71560;
	#10 counter$count = 71561;
	#10 counter$count = 71562;
	#10 counter$count = 71563;
	#10 counter$count = 71564;
	#10 counter$count = 71565;
	#10 counter$count = 71566;
	#10 counter$count = 71567;
	#10 counter$count = 71568;
	#10 counter$count = 71569;
	#10 counter$count = 71570;
	#10 counter$count = 71571;
	#10 counter$count = 71572;
	#10 counter$count = 71573;
	#10 counter$count = 71574;
	#10 counter$count = 71575;
	#10 counter$count = 71576;
	#10 counter$count = 71577;
	#10 counter$count = 71578;
	#10 counter$count = 71579;
	#10 counter$count = 71580;
	#10 counter$count = 71581;
	#10 counter$count = 71582;
	#10 counter$count = 71583;
	#10 counter$count = 71584;
	#10 counter$count = 71585;
	#10 counter$count = 71586;
	#10 counter$count = 71587;
	#10 counter$count = 71588;
	#10 counter$count = 71589;
	#10 counter$count = 71590;
	#10 counter$count = 71591;
	#10 counter$count = 71592;
	#10 counter$count = 71593;
	#10 counter$count = 71594;
	#10 counter$count = 71595;
	#10 counter$count = 71596;
	#10 counter$count = 71597;
	#10 counter$count = 71598;
	#10 counter$count = 71599;
	#10 counter$count = 71600;
	#10 counter$count = 71601;
	#10 counter$count = 71602;
	#10 counter$count = 71603;
	#10 counter$count = 71604;
	#10 counter$count = 71605;
	#10 counter$count = 71606;
	#10 counter$count = 71607;
	#10 counter$count = 71608;
	#10 counter$count = 71609;
	#10 counter$count = 71610;
	#10 counter$count = 71611;
	#10 counter$count = 71612;
	#10 counter$count = 71613;
	#10 counter$count = 71614;
	#10 counter$count = 71615;
	#10 counter$count = 71616;
	#10 counter$count = 71617;
	#10 counter$count = 71618;
	#10 counter$count = 71619;
	#10 counter$count = 71620;
	#10 counter$count = 71621;
	#10 counter$count = 71622;
	#10 counter$count = 71623;
	#10 counter$count = 71624;
	#10 counter$count = 71625;
	#10 counter$count = 71626;
	#10 counter$count = 71627;
	#10 counter$count = 71628;
	#10 counter$count = 71629;
	#10 counter$count = 71630;
	#10 counter$count = 71631;
	#10 counter$count = 71632;
	#10 counter$count = 71633;
	#10 counter$count = 71634;
	#10 counter$count = 71635;
	#10 counter$count = 71636;
	#10 counter$count = 71637;
	#10 counter$count = 71638;
	#10 counter$count = 71639;
	#10 counter$count = 71640;
	#10 counter$count = 71641;
	#10 counter$count = 71642;
	#10 counter$count = 71643;
	#10 counter$count = 71644;
	#10 counter$count = 71645;
	#10 counter$count = 71646;
	#10 counter$count = 71647;
	#10 counter$count = 71648;
	#10 counter$count = 71649;
	#10 counter$count = 71650;
	#10 counter$count = 71651;
	#10 counter$count = 71652;
	#10 counter$count = 71653;
	#10 counter$count = 71654;
	#10 counter$count = 71655;
	#10 counter$count = 71656;
	#10 counter$count = 71657;
	#10 counter$count = 71658;
	#10 counter$count = 71659;
	#10 counter$count = 71660;
	#10 counter$count = 71661;
	#10 counter$count = 71662;
	#10 counter$count = 71663;
	#10 counter$count = 71664;
	#10 counter$count = 71665;
	#10 counter$count = 71666;
	#10 counter$count = 71667;
	#10 counter$count = 71668;
	#10 counter$count = 71669;
	#10 counter$count = 71670;
	#10 counter$count = 71671;
	#10 counter$count = 71672;
	#10 counter$count = 71673;
	#10 counter$count = 71674;
	#10 counter$count = 71675;
	#10 counter$count = 71676;
	#10 counter$count = 71677;
	#10 counter$count = 71678;
	#10 counter$count = 71679;
	#10 counter$count = 71680;
	#10 counter$count = 71681;
	#10 counter$count = 71682;
	#10 counter$count = 71683;
	#10 counter$count = 71684;
	#10 counter$count = 71685;
	#10 counter$count = 71686;
	#10 counter$count = 71687;
	#10 counter$count = 71688;
	#10 counter$count = 71689;
	#10 counter$count = 71690;
	#10 counter$count = 71691;
	#10 counter$count = 71692;
	#10 counter$count = 71693;
	#10 counter$count = 71694;
	#10 counter$count = 71695;
	#10 counter$count = 71696;
	#10 counter$count = 71697;
	#10 counter$count = 71698;
	#10 counter$count = 71699;
	#10 counter$count = 71700;
	#10 counter$count = 71701;
	#10 counter$count = 71702;
	#10 counter$count = 71703;
	#10 counter$count = 71704;
	#10 counter$count = 71705;
	#10 counter$count = 71706;
	#10 counter$count = 71707;
	#10 counter$count = 71708;
	#10 counter$count = 71709;
	#10 counter$count = 71710;
	#10 counter$count = 71711;
	#10 counter$count = 71712;
	#10 counter$count = 71713;
	#10 counter$count = 71714;
	#10 counter$count = 71715;
	#10 counter$count = 71716;
	#10 counter$count = 71717;
	#10 counter$count = 71718;
	#10 counter$count = 71719;
	#10 counter$count = 71720;
	#10 counter$count = 71721;
	#10 counter$count = 71722;
	#10 counter$count = 71723;
	#10 counter$count = 71724;
	#10 counter$count = 71725;
	#10 counter$count = 71726;
	#10 counter$count = 71727;
	#10 counter$count = 71728;
	#10 counter$count = 71729;
	#10 counter$count = 71730;
	#10 counter$count = 71731;
	#10 counter$count = 71732;
	#10 counter$count = 71733;
	#10 counter$count = 71734;
	#10 counter$count = 71735;
	#10 counter$count = 71736;
	#10 counter$count = 71737;
	#10 counter$count = 71738;
	#10 counter$count = 71739;
	#10 counter$count = 71740;
	#10 counter$count = 71741;
	#10 counter$count = 71742;
	#10 counter$count = 71743;
	#10 counter$count = 71744;
	#10 counter$count = 71745;
	#10 counter$count = 71746;
	#10 counter$count = 71747;
	#10 counter$count = 71748;
	#10 counter$count = 71749;
	#10 counter$count = 71750;
	#10 counter$count = 71751;
	#10 counter$count = 71752;
	#10 counter$count = 71753;
	#10 counter$count = 71754;
	#10 counter$count = 71755;
	#10 counter$count = 71756;
	#10 counter$count = 71757;
	#10 counter$count = 71758;
	#10 counter$count = 71759;
	#10 counter$count = 71760;
	#10 counter$count = 71761;
	#10 counter$count = 71762;
	#10 counter$count = 71763;
	#10 counter$count = 71764;
	#10 counter$count = 71765;
	#10 counter$count = 71766;
	#10 counter$count = 71767;
	#10 counter$count = 71768;
	#10 counter$count = 71769;
	#10 counter$count = 71770;
	#10 counter$count = 71771;
	#10 counter$count = 71772;
	#10 counter$count = 71773;
	#10 counter$count = 71774;
	#10 counter$count = 71775;
	#10 counter$count = 71776;
	#10 counter$count = 71777;
	#10 counter$count = 71778;
	#10 counter$count = 71779;
	#10 counter$count = 71780;
	#10 counter$count = 71781;
	#10 counter$count = 71782;
	#10 counter$count = 71783;
	#10 counter$count = 71784;
	#10 counter$count = 71785;
	#10 counter$count = 71786;
	#10 counter$count = 71787;
	#10 counter$count = 71788;
	#10 counter$count = 71789;
	#10 counter$count = 71790;
	#10 counter$count = 71791;
	#10 counter$count = 71792;
	#10 counter$count = 71793;
	#10 counter$count = 71794;
	#10 counter$count = 71795;
	#10 counter$count = 71796;
	#10 counter$count = 71797;
	#10 counter$count = 71798;
	#10 counter$count = 71799;
	#10 counter$count = 71800;
	#10 counter$count = 71801;
	#10 counter$count = 71802;
	#10 counter$count = 71803;
	#10 counter$count = 71804;
	#10 counter$count = 71805;
	#10 counter$count = 71806;
	#10 counter$count = 71807;
	#10 counter$count = 71808;
	#10 counter$count = 71809;
	#10 counter$count = 71810;
	#10 counter$count = 71811;
	#10 counter$count = 71812;
	#10 counter$count = 71813;
	#10 counter$count = 71814;
	#10 counter$count = 71815;
	#10 counter$count = 71816;
	#10 counter$count = 71817;
	#10 counter$count = 71818;
	#10 counter$count = 71819;
	#10 counter$count = 71820;
	#10 counter$count = 71821;
	#10 counter$count = 71822;
	#10 counter$count = 71823;
	#10 counter$count = 71824;
	#10 counter$count = 71825;
	#10 counter$count = 71826;
	#10 counter$count = 71827;
	#10 counter$count = 71828;
	#10 counter$count = 71829;
	#10 counter$count = 71830;
	#10 counter$count = 71831;
	#10 counter$count = 71832;
	#10 counter$count = 71833;
	#10 counter$count = 71834;
	#10 counter$count = 71835;
	#10 counter$count = 71836;
	#10 counter$count = 71837;
	#10 counter$count = 71838;
	#10 counter$count = 71839;
	#10 counter$count = 71840;
	#10 counter$count = 71841;
	#10 counter$count = 71842;
	#10 counter$count = 71843;
	#10 counter$count = 71844;
	#10 counter$count = 71845;
	#10 counter$count = 71846;
	#10 counter$count = 71847;
	#10 counter$count = 71848;
	#10 counter$count = 71849;
	#10 counter$count = 71850;
	#10 counter$count = 71851;
	#10 counter$count = 71852;
	#10 counter$count = 71853;
	#10 counter$count = 71854;
	#10 counter$count = 71855;
	#10 counter$count = 71856;
	#10 counter$count = 71857;
	#10 counter$count = 71858;
	#10 counter$count = 71859;
	#10 counter$count = 71860;
	#10 counter$count = 71861;
	#10 counter$count = 71862;
	#10 counter$count = 71863;
	#10 counter$count = 71864;
	#10 counter$count = 71865;
	#10 counter$count = 71866;
	#10 counter$count = 71867;
	#10 counter$count = 71868;
	#10 counter$count = 71869;
	#10 counter$count = 71870;
	#10 counter$count = 71871;
	#10 counter$count = 71872;
	#10 counter$count = 71873;
	#10 counter$count = 71874;
	#10 counter$count = 71875;
	#10 counter$count = 71876;
	#10 counter$count = 71877;
	#10 counter$count = 71878;
	#10 counter$count = 71879;
	#10 counter$count = 71880;
	#10 counter$count = 71881;
	#10 counter$count = 71882;
	#10 counter$count = 71883;
	#10 counter$count = 71884;
	#10 counter$count = 71885;
	#10 counter$count = 71886;
	#10 counter$count = 71887;
	#10 counter$count = 71888;
	#10 counter$count = 71889;
	#10 counter$count = 71890;
	#10 counter$count = 71891;
	#10 counter$count = 71892;
	#10 counter$count = 71893;
	#10 counter$count = 71894;
	#10 counter$count = 71895;
	#10 counter$count = 71896;
	#10 counter$count = 71897;
	#10 counter$count = 71898;
	#10 counter$count = 71899;
	#10 counter$count = 71900;
	#10 counter$count = 71901;
	#10 counter$count = 71902;
	#10 counter$count = 71903;
	#10 counter$count = 71904;
	#10 counter$count = 71905;
	#10 counter$count = 71906;
	#10 counter$count = 71907;
	#10 counter$count = 71908;
	#10 counter$count = 71909;
	#10 counter$count = 71910;
	#10 counter$count = 71911;
	#10 counter$count = 71912;
	#10 counter$count = 71913;
	#10 counter$count = 71914;
	#10 counter$count = 71915;
	#10 counter$count = 71916;
	#10 counter$count = 71917;
	#10 counter$count = 71918;
	#10 counter$count = 71919;
	#10 counter$count = 71920;
	#10 counter$count = 71921;
	#10 counter$count = 71922;
	#10 counter$count = 71923;
	#10 counter$count = 71924;
	#10 counter$count = 71925;
	#10 counter$count = 71926;
	#10 counter$count = 71927;
	#10 counter$count = 71928;
	#10 counter$count = 71929;
	#10 counter$count = 71930;
	#10 counter$count = 71931;
	#10 counter$count = 71932;
	#10 counter$count = 71933;
	#10 counter$count = 71934;
	#10 counter$count = 71935;
	#10 counter$count = 71936;
	#10 counter$count = 71937;
	#10 counter$count = 71938;
	#10 counter$count = 71939;
	#10 counter$count = 71940;
	#10 counter$count = 71941;
	#10 counter$count = 71942;
	#10 counter$count = 71943;
	#10 counter$count = 71944;
	#10 counter$count = 71945;
	#10 counter$count = 71946;
	#10 counter$count = 71947;
	#10 counter$count = 71948;
	#10 counter$count = 71949;
	#10 counter$count = 71950;
	#10 counter$count = 71951;
	#10 counter$count = 71952;
	#10 counter$count = 71953;
	#10 counter$count = 71954;
	#10 counter$count = 71955;
	#10 counter$count = 71956;
	#10 counter$count = 71957;
	#10 counter$count = 71958;
	#10 counter$count = 71959;
	#10 counter$count = 71960;
	#10 counter$count = 71961;
	#10 counter$count = 71962;
	#10 counter$count = 71963;
	#10 counter$count = 71964;
	#10 counter$count = 71965;
	#10 counter$count = 71966;
	#10 counter$count = 71967;
	#10 counter$count = 71968;
	#10 counter$count = 71969;
	#10 counter$count = 71970;
	#10 counter$count = 71971;
	#10 counter$count = 71972;
	#10 counter$count = 71973;
	#10 counter$count = 71974;
	#10 counter$count = 71975;
	#10 counter$count = 71976;
	#10 counter$count = 71977;
	#10 counter$count = 71978;
	#10 counter$count = 71979;
	#10 counter$count = 71980;
	#10 counter$count = 71981;
	#10 counter$count = 71982;
	#10 counter$count = 71983;
	#10 counter$count = 71984;
	#10 counter$count = 71985;
	#10 counter$count = 71986;
	#10 counter$count = 71987;
	#10 counter$count = 71988;
	#10 counter$count = 71989;
	#10 counter$count = 71990;
	#10 counter$count = 71991;
	#10 counter$count = 71992;
	#10 counter$count = 71993;
	#10 counter$count = 71994;
	#10 counter$count = 71995;
	#10 counter$count = 71996;
	#10 counter$count = 71997;
	#10 counter$count = 71998;
	#10 counter$count = 71999;
	#10 counter$count = 72000;
	#10 counter$count = 72001;
	#10 counter$count = 72002;
	#10 counter$count = 72003;
	#10 counter$count = 72004;
	#10 counter$count = 72005;
	#10 counter$count = 72006;
	#10 counter$count = 72007;
	#10 counter$count = 72008;
	#10 counter$count = 72009;
	#10 counter$count = 72010;
	#10 counter$count = 72011;
	#10 counter$count = 72012;
	#10 counter$count = 72013;
	#10 counter$count = 72014;
	#10 counter$count = 72015;
	#10 counter$count = 72016;
	#10 counter$count = 72017;
	#10 counter$count = 72018;
	#10 counter$count = 72019;
	#10 counter$count = 72020;
	#10 counter$count = 72021;
	#10 counter$count = 72022;
	#10 counter$count = 72023;
	#10 counter$count = 72024;
	#10 counter$count = 72025;
	#10 counter$count = 72026;
	#10 counter$count = 72027;
	#10 counter$count = 72028;
	#10 counter$count = 72029;
	#10 counter$count = 72030;
	#10 counter$count = 72031;
	#10 counter$count = 72032;
	#10 counter$count = 72033;
	#10 counter$count = 72034;
	#10 counter$count = 72035;
	#10 counter$count = 72036;
	#10 counter$count = 72037;
	#10 counter$count = 72038;
	#10 counter$count = 72039;
	#10 counter$count = 72040;
	#10 counter$count = 72041;
	#10 counter$count = 72042;
	#10 counter$count = 72043;
	#10 counter$count = 72044;
	#10 counter$count = 72045;
	#10 counter$count = 72046;
	#10 counter$count = 72047;
	#10 counter$count = 72048;
	#10 counter$count = 72049;
	#10 counter$count = 72050;
	#10 counter$count = 72051;
	#10 counter$count = 72052;
	#10 counter$count = 72053;
	#10 counter$count = 72054;
	#10 counter$count = 72055;
	#10 counter$count = 72056;
	#10 counter$count = 72057;
	#10 counter$count = 72058;
	#10 counter$count = 72059;
	#10 counter$count = 72060;
	#10 counter$count = 72061;
	#10 counter$count = 72062;
	#10 counter$count = 72063;
	#10 counter$count = 72064;
	#10 counter$count = 72065;
	#10 counter$count = 72066;
	#10 counter$count = 72067;
	#10 counter$count = 72068;
	#10 counter$count = 72069;
	#10 counter$count = 72070;
	#10 counter$count = 72071;
	#10 counter$count = 72072;
	#10 counter$count = 72073;
	#10 counter$count = 72074;
	#10 counter$count = 72075;
	#10 counter$count = 72076;
	#10 counter$count = 72077;
	#10 counter$count = 72078;
	#10 counter$count = 72079;
	#10 counter$count = 72080;
	#10 counter$count = 72081;
	#10 counter$count = 72082;
	#10 counter$count = 72083;
	#10 counter$count = 72084;
	#10 counter$count = 72085;
	#10 counter$count = 72086;
	#10 counter$count = 72087;
	#10 counter$count = 72088;
	#10 counter$count = 72089;
	#10 counter$count = 72090;
	#10 counter$count = 72091;
	#10 counter$count = 72092;
	#10 counter$count = 72093;
	#10 counter$count = 72094;
	#10 counter$count = 72095;
	#10 counter$count = 72096;
	#10 counter$count = 72097;
	#10 counter$count = 72098;
	#10 counter$count = 72099;
	#10 counter$count = 72100;
	#10 counter$count = 72101;
	#10 counter$count = 72102;
	#10 counter$count = 72103;
	#10 counter$count = 72104;
	#10 counter$count = 72105;
	#10 counter$count = 72106;
	#10 counter$count = 72107;
	#10 counter$count = 72108;
	#10 counter$count = 72109;
	#10 counter$count = 72110;
	#10 counter$count = 72111;
	#10 counter$count = 72112;
	#10 counter$count = 72113;
	#10 counter$count = 72114;
	#10 counter$count = 72115;
	#10 counter$count = 72116;
	#10 counter$count = 72117;
	#10 counter$count = 72118;
	#10 counter$count = 72119;
	#10 counter$count = 72120;
	#10 counter$count = 72121;
	#10 counter$count = 72122;
	#10 counter$count = 72123;
	#10 counter$count = 72124;
	#10 counter$count = 72125;
	#10 counter$count = 72126;
	#10 counter$count = 72127;
	#10 counter$count = 72128;
	#10 counter$count = 72129;
	#10 counter$count = 72130;
	#10 counter$count = 72131;
	#10 counter$count = 72132;
	#10 counter$count = 72133;
	#10 counter$count = 72134;
	#10 counter$count = 72135;
	#10 counter$count = 72136;
	#10 counter$count = 72137;
	#10 counter$count = 72138;
	#10 counter$count = 72139;
	#10 counter$count = 72140;
	#10 counter$count = 72141;
	#10 counter$count = 72142;
	#10 counter$count = 72143;
	#10 counter$count = 72144;
	#10 counter$count = 72145;
	#10 counter$count = 72146;
	#10 counter$count = 72147;
	#10 counter$count = 72148;
	#10 counter$count = 72149;
	#10 counter$count = 72150;
	#10 counter$count = 72151;
	#10 counter$count = 72152;
	#10 counter$count = 72153;
	#10 counter$count = 72154;
	#10 counter$count = 72155;
	#10 counter$count = 72156;
	#10 counter$count = 72157;
	#10 counter$count = 72158;
	#10 counter$count = 72159;
	#10 counter$count = 72160;
	#10 counter$count = 72161;
	#10 counter$count = 72162;
	#10 counter$count = 72163;
	#10 counter$count = 72164;
	#10 counter$count = 72165;
	#10 counter$count = 72166;
	#10 counter$count = 72167;
	#10 counter$count = 72168;
	#10 counter$count = 72169;
	#10 counter$count = 72170;
	#10 counter$count = 72171;
	#10 counter$count = 72172;
	#10 counter$count = 72173;
	#10 counter$count = 72174;
	#10 counter$count = 72175;
	#10 counter$count = 72176;
	#10 counter$count = 72177;
	#10 counter$count = 72178;
	#10 counter$count = 72179;
	#10 counter$count = 72180;
	#10 counter$count = 72181;
	#10 counter$count = 72182;
	#10 counter$count = 72183;
	#10 counter$count = 72184;
	#10 counter$count = 72185;
	#10 counter$count = 72186;
	#10 counter$count = 72187;
	#10 counter$count = 72188;
	#10 counter$count = 72189;
	#10 counter$count = 72190;
	#10 counter$count = 72191;
	#10 counter$count = 72192;
	#10 counter$count = 72193;
	#10 counter$count = 72194;
	#10 counter$count = 72195;
	#10 counter$count = 72196;
	#10 counter$count = 72197;
	#10 counter$count = 72198;
	#10 counter$count = 72199;
	#10 counter$count = 72200;
	#10 counter$count = 72201;
	#10 counter$count = 72202;
	#10 counter$count = 72203;
	#10 counter$count = 72204;
	#10 counter$count = 72205;
	#10 counter$count = 72206;
	#10 counter$count = 72207;
	#10 counter$count = 72208;
	#10 counter$count = 72209;
	#10 counter$count = 72210;
	#10 counter$count = 72211;
	#10 counter$count = 72212;
	#10 counter$count = 72213;
	#10 counter$count = 72214;
	#10 counter$count = 72215;
	#10 counter$count = 72216;
	#10 counter$count = 72217;
	#10 counter$count = 72218;
	#10 counter$count = 72219;
	#10 counter$count = 72220;
	#10 counter$count = 72221;
	#10 counter$count = 72222;
	#10 counter$count = 72223;
	#10 counter$count = 72224;
	#10 counter$count = 72225;
	#10 counter$count = 72226;
	#10 counter$count = 72227;
	#10 counter$count = 72228;
	#10 counter$count = 72229;
	#10 counter$count = 72230;
	#10 counter$count = 72231;
	#10 counter$count = 72232;
	#10 counter$count = 72233;
	#10 counter$count = 72234;
	#10 counter$count = 72235;
	#10 counter$count = 72236;
	#10 counter$count = 72237;
	#10 counter$count = 72238;
	#10 counter$count = 72239;
	#10 counter$count = 72240;
	#10 counter$count = 72241;
	#10 counter$count = 72242;
	#10 counter$count = 72243;
	#10 counter$count = 72244;
	#10 counter$count = 72245;
	#10 counter$count = 72246;
	#10 counter$count = 72247;
	#10 counter$count = 72248;
	#10 counter$count = 72249;
	#10 counter$count = 72250;
	#10 counter$count = 72251;
	#10 counter$count = 72252;
	#10 counter$count = 72253;
	#10 counter$count = 72254;
	#10 counter$count = 72255;
	#10 counter$count = 72256;
	#10 counter$count = 72257;
	#10 counter$count = 72258;
	#10 counter$count = 72259;
	#10 counter$count = 72260;
	#10 counter$count = 72261;
	#10 counter$count = 72262;
	#10 counter$count = 72263;
	#10 counter$count = 72264;
	#10 counter$count = 72265;
	#10 counter$count = 72266;
	#10 counter$count = 72267;
	#10 counter$count = 72268;
	#10 counter$count = 72269;
	#10 counter$count = 72270;
	#10 counter$count = 72271;
	#10 counter$count = 72272;
	#10 counter$count = 72273;
	#10 counter$count = 72274;
	#10 counter$count = 72275;
	#10 counter$count = 72276;
	#10 counter$count = 72277;
	#10 counter$count = 72278;
	#10 counter$count = 72279;
	#10 counter$count = 72280;
	#10 counter$count = 72281;
	#10 counter$count = 72282;
	#10 counter$count = 72283;
	#10 counter$count = 72284;
	#10 counter$count = 72285;
	#10 counter$count = 72286;
	#10 counter$count = 72287;
	#10 counter$count = 72288;
	#10 counter$count = 72289;
	#10 counter$count = 72290;
	#10 counter$count = 72291;
	#10 counter$count = 72292;
	#10 counter$count = 72293;
	#10 counter$count = 72294;
	#10 counter$count = 72295;
	#10 counter$count = 72296;
	#10 counter$count = 72297;
	#10 counter$count = 72298;
	#10 counter$count = 72299;
	#10 counter$count = 72300;
	#10 counter$count = 72301;
	#10 counter$count = 72302;
	#10 counter$count = 72303;
	#10 counter$count = 72304;
	#10 counter$count = 72305;
	#10 counter$count = 72306;
	#10 counter$count = 72307;
	#10 counter$count = 72308;
	#10 counter$count = 72309;
	#10 counter$count = 72310;
	#10 counter$count = 72311;
	#10 counter$count = 72312;
	#10 counter$count = 72313;
	#10 counter$count = 72314;
	#10 counter$count = 72315;
	#10 counter$count = 72316;
	#10 counter$count = 72317;
	#10 counter$count = 72318;
	#10 counter$count = 72319;
	#10 counter$count = 72320;
	#10 counter$count = 72321;
	#10 counter$count = 72322;
	#10 counter$count = 72323;
	#10 counter$count = 72324;
	#10 counter$count = 72325;
	#10 counter$count = 72326;
	#10 counter$count = 72327;
	#10 counter$count = 72328;
	#10 counter$count = 72329;
	#10 counter$count = 72330;
	#10 counter$count = 72331;
	#10 counter$count = 72332;
	#10 counter$count = 72333;
	#10 counter$count = 72334;
	#10 counter$count = 72335;
	#10 counter$count = 72336;
	#10 counter$count = 72337;
	#10 counter$count = 72338;
	#10 counter$count = 72339;
	#10 counter$count = 72340;
	#10 counter$count = 72341;
	#10 counter$count = 72342;
	#10 counter$count = 72343;
	#10 counter$count = 72344;
	#10 counter$count = 72345;
	#10 counter$count = 72346;
	#10 counter$count = 72347;
	#10 counter$count = 72348;
	#10 counter$count = 72349;
	#10 counter$count = 72350;
	#10 counter$count = 72351;
	#10 counter$count = 72352;
	#10 counter$count = 72353;
	#10 counter$count = 72354;
	#10 counter$count = 72355;
	#10 counter$count = 72356;
	#10 counter$count = 72357;
	#10 counter$count = 72358;
	#10 counter$count = 72359;
	#10 counter$count = 72360;
	#10 counter$count = 72361;
	#10 counter$count = 72362;
	#10 counter$count = 72363;
	#10 counter$count = 72364;
	#10 counter$count = 72365;
	#10 counter$count = 72366;
	#10 counter$count = 72367;
	#10 counter$count = 72368;
	#10 counter$count = 72369;
	#10 counter$count = 72370;
	#10 counter$count = 72371;
	#10 counter$count = 72372;
	#10 counter$count = 72373;
	#10 counter$count = 72374;
	#10 counter$count = 72375;
	#10 counter$count = 72376;
	#10 counter$count = 72377;
	#10 counter$count = 72378;
	#10 counter$count = 72379;
	#10 counter$count = 72380;
	#10 counter$count = 72381;
	#10 counter$count = 72382;
	#10 counter$count = 72383;
	#10 counter$count = 72384;
	#10 counter$count = 72385;
	#10 counter$count = 72386;
	#10 counter$count = 72387;
	#10 counter$count = 72388;
	#10 counter$count = 72389;
	#10 counter$count = 72390;
	#10 counter$count = 72391;
	#10 counter$count = 72392;
	#10 counter$count = 72393;
	#10 counter$count = 72394;
	#10 counter$count = 72395;
	#10 counter$count = 72396;
	#10 counter$count = 72397;
	#10 counter$count = 72398;
	#10 counter$count = 72399;
	#10 counter$count = 72400;
	#10 counter$count = 72401;
	#10 counter$count = 72402;
	#10 counter$count = 72403;
	#10 counter$count = 72404;
	#10 counter$count = 72405;
	#10 counter$count = 72406;
	#10 counter$count = 72407;
	#10 counter$count = 72408;
	#10 counter$count = 72409;
	#10 counter$count = 72410;
	#10 counter$count = 72411;
	#10 counter$count = 72412;
	#10 counter$count = 72413;
	#10 counter$count = 72414;
	#10 counter$count = 72415;
	#10 counter$count = 72416;
	#10 counter$count = 72417;
	#10 counter$count = 72418;
	#10 counter$count = 72419;
	#10 counter$count = 72420;
	#10 counter$count = 72421;
	#10 counter$count = 72422;
	#10 counter$count = 72423;
	#10 counter$count = 72424;
	#10 counter$count = 72425;
	#10 counter$count = 72426;
	#10 counter$count = 72427;
	#10 counter$count = 72428;
	#10 counter$count = 72429;
	#10 counter$count = 72430;
	#10 counter$count = 72431;
	#10 counter$count = 72432;
	#10 counter$count = 72433;
	#10 counter$count = 72434;
	#10 counter$count = 72435;
	#10 counter$count = 72436;
	#10 counter$count = 72437;
	#10 counter$count = 72438;
	#10 counter$count = 72439;
	#10 counter$count = 72440;
	#10 counter$count = 72441;
	#10 counter$count = 72442;
	#10 counter$count = 72443;
	#10 counter$count = 72444;
	#10 counter$count = 72445;
	#10 counter$count = 72446;
	#10 counter$count = 72447;
	#10 counter$count = 72448;
	#10 counter$count = 72449;
	#10 counter$count = 72450;
	#10 counter$count = 72451;
	#10 counter$count = 72452;
	#10 counter$count = 72453;
	#10 counter$count = 72454;
	#10 counter$count = 72455;
	#10 counter$count = 72456;
	#10 counter$count = 72457;
	#10 counter$count = 72458;
	#10 counter$count = 72459;
	#10 counter$count = 72460;
	#10 counter$count = 72461;
	#10 counter$count = 72462;
	#10 counter$count = 72463;
	#10 counter$count = 72464;
	#10 counter$count = 72465;
	#10 counter$count = 72466;
	#10 counter$count = 72467;
	#10 counter$count = 72468;
	#10 counter$count = 72469;
	#10 counter$count = 72470;
	#10 counter$count = 72471;
	#10 counter$count = 72472;
	#10 counter$count = 72473;
	#10 counter$count = 72474;
	#10 counter$count = 72475;
	#10 counter$count = 72476;
	#10 counter$count = 72477;
	#10 counter$count = 72478;
	#10 counter$count = 72479;
	#10 counter$count = 72480;
	#10 counter$count = 72481;
	#10 counter$count = 72482;
	#10 counter$count = 72483;
	#10 counter$count = 72484;
	#10 counter$count = 72485;
	#10 counter$count = 72486;
	#10 counter$count = 72487;
	#10 counter$count = 72488;
	#10 counter$count = 72489;
	#10 counter$count = 72490;
	#10 counter$count = 72491;
	#10 counter$count = 72492;
	#10 counter$count = 72493;
	#10 counter$count = 72494;
	#10 counter$count = 72495;
	#10 counter$count = 72496;
	#10 counter$count = 72497;
	#10 counter$count = 72498;
	#10 counter$count = 72499;
	#10 counter$count = 72500;
	#10 counter$count = 72501;
	#10 counter$count = 72502;
	#10 counter$count = 72503;
	#10 counter$count = 72504;
	#10 counter$count = 72505;
	#10 counter$count = 72506;
	#10 counter$count = 72507;
	#10 counter$count = 72508;
	#10 counter$count = 72509;
	#10 counter$count = 72510;
	#10 counter$count = 72511;
	#10 counter$count = 72512;
	#10 counter$count = 72513;
	#10 counter$count = 72514;
	#10 counter$count = 72515;
	#10 counter$count = 72516;
	#10 counter$count = 72517;
	#10 counter$count = 72518;
	#10 counter$count = 72519;
	#10 counter$count = 72520;
	#10 counter$count = 72521;
	#10 counter$count = 72522;
	#10 counter$count = 72523;
	#10 counter$count = 72524;
	#10 counter$count = 72525;
	#10 counter$count = 72526;
	#10 counter$count = 72527;
	#10 counter$count = 72528;
	#10 counter$count = 72529;
	#10 counter$count = 72530;
	#10 counter$count = 72531;
	#10 counter$count = 72532;
	#10 counter$count = 72533;
	#10 counter$count = 72534;
	#10 counter$count = 72535;
	#10 counter$count = 72536;
	#10 counter$count = 72537;
	#10 counter$count = 72538;
	#10 counter$count = 72539;
	#10 counter$count = 72540;
	#10 counter$count = 72541;
	#10 counter$count = 72542;
	#10 counter$count = 72543;
	#10 counter$count = 72544;
	#10 counter$count = 72545;
	#10 counter$count = 72546;
	#10 counter$count = 72547;
	#10 counter$count = 72548;
	#10 counter$count = 72549;
	#10 counter$count = 72550;
	#10 counter$count = 72551;
	#10 counter$count = 72552;
	#10 counter$count = 72553;
	#10 counter$count = 72554;
	#10 counter$count = 72555;
	#10 counter$count = 72556;
	#10 counter$count = 72557;
	#10 counter$count = 72558;
	#10 counter$count = 72559;
	#10 counter$count = 72560;
	#10 counter$count = 72561;
	#10 counter$count = 72562;
	#10 counter$count = 72563;
	#10 counter$count = 72564;
	#10 counter$count = 72565;
	#10 counter$count = 72566;
	#10 counter$count = 72567;
	#10 counter$count = 72568;
	#10 counter$count = 72569;
	#10 counter$count = 72570;
	#10 counter$count = 72571;
	#10 counter$count = 72572;
	#10 counter$count = 72573;
	#10 counter$count = 72574;
	#10 counter$count = 72575;
	#10 counter$count = 72576;
	#10 counter$count = 72577;
	#10 counter$count = 72578;
	#10 counter$count = 72579;
	#10 counter$count = 72580;
	#10 counter$count = 72581;
	#10 counter$count = 72582;
	#10 counter$count = 72583;
	#10 counter$count = 72584;
	#10 counter$count = 72585;
	#10 counter$count = 72586;
	#10 counter$count = 72587;
	#10 counter$count = 72588;
	#10 counter$count = 72589;
	#10 counter$count = 72590;
	#10 counter$count = 72591;
	#10 counter$count = 72592;
	#10 counter$count = 72593;
	#10 counter$count = 72594;
	#10 counter$count = 72595;
	#10 counter$count = 72596;
	#10 counter$count = 72597;
	#10 counter$count = 72598;
	#10 counter$count = 72599;
	#10 counter$count = 72600;
	#10 counter$count = 72601;
	#10 counter$count = 72602;
	#10 counter$count = 72603;
	#10 counter$count = 72604;
	#10 counter$count = 72605;
	#10 counter$count = 72606;
	#10 counter$count = 72607;
	#10 counter$count = 72608;
	#10 counter$count = 72609;
	#10 counter$count = 72610;
	#10 counter$count = 72611;
	#10 counter$count = 72612;
	#10 counter$count = 72613;
	#10 counter$count = 72614;
	#10 counter$count = 72615;
	#10 counter$count = 72616;
	#10 counter$count = 72617;
	#10 counter$count = 72618;
	#10 counter$count = 72619;
	#10 counter$count = 72620;
	#10 counter$count = 72621;
	#10 counter$count = 72622;
	#10 counter$count = 72623;
	#10 counter$count = 72624;
	#10 counter$count = 72625;
	#10 counter$count = 72626;
	#10 counter$count = 72627;
	#10 counter$count = 72628;
	#10 counter$count = 72629;
	#10 counter$count = 72630;
	#10 counter$count = 72631;
	#10 counter$count = 72632;
	#10 counter$count = 72633;
	#10 counter$count = 72634;
	#10 counter$count = 72635;
	#10 counter$count = 72636;
	#10 counter$count = 72637;
	#10 counter$count = 72638;
	#10 counter$count = 72639;
	#10 counter$count = 72640;
	#10 counter$count = 72641;
	#10 counter$count = 72642;
	#10 counter$count = 72643;
	#10 counter$count = 72644;
	#10 counter$count = 72645;
	#10 counter$count = 72646;
	#10 counter$count = 72647;
	#10 counter$count = 72648;
	#10 counter$count = 72649;
	#10 counter$count = 72650;
	#10 counter$count = 72651;
	#10 counter$count = 72652;
	#10 counter$count = 72653;
	#10 counter$count = 72654;
	#10 counter$count = 72655;
	#10 counter$count = 72656;
	#10 counter$count = 72657;
	#10 counter$count = 72658;
	#10 counter$count = 72659;
	#10 counter$count = 72660;
	#10 counter$count = 72661;
	#10 counter$count = 72662;
	#10 counter$count = 72663;
	#10 counter$count = 72664;
	#10 counter$count = 72665;
	#10 counter$count = 72666;
	#10 counter$count = 72667;
	#10 counter$count = 72668;
	#10 counter$count = 72669;
	#10 counter$count = 72670;
	#10 counter$count = 72671;
	#10 counter$count = 72672;
	#10 counter$count = 72673;
	#10 counter$count = 72674;
	#10 counter$count = 72675;
	#10 counter$count = 72676;
	#10 counter$count = 72677;
	#10 counter$count = 72678;
	#10 counter$count = 72679;
	#10 counter$count = 72680;
	#10 counter$count = 72681;
	#10 counter$count = 72682;
	#10 counter$count = 72683;
	#10 counter$count = 72684;
	#10 counter$count = 72685;
	#10 counter$count = 72686;
	#10 counter$count = 72687;
	#10 counter$count = 72688;
	#10 counter$count = 72689;
	#10 counter$count = 72690;
	#10 counter$count = 72691;
	#10 counter$count = 72692;
	#10 counter$count = 72693;
	#10 counter$count = 72694;
	#10 counter$count = 72695;
	#10 counter$count = 72696;
	#10 counter$count = 72697;
	#10 counter$count = 72698;
	#10 counter$count = 72699;
	#10 counter$count = 72700;
	#10 counter$count = 72701;
	#10 counter$count = 72702;
	#10 counter$count = 72703;
	#10 counter$count = 72704;
	#10 counter$count = 72705;
	#10 counter$count = 72706;
	#10 counter$count = 72707;
	#10 counter$count = 72708;
	#10 counter$count = 72709;
	#10 counter$count = 72710;
	#10 counter$count = 72711;
	#10 counter$count = 72712;
	#10 counter$count = 72713;
	#10 counter$count = 72714;
	#10 counter$count = 72715;
	#10 counter$count = 72716;
	#10 counter$count = 72717;
	#10 counter$count = 72718;
	#10 counter$count = 72719;
	#10 counter$count = 72720;
	#10 counter$count = 72721;
	#10 counter$count = 72722;
	#10 counter$count = 72723;
	#10 counter$count = 72724;
	#10 counter$count = 72725;
	#10 counter$count = 72726;
	#10 counter$count = 72727;
	#10 counter$count = 72728;
	#10 counter$count = 72729;
	#10 counter$count = 72730;
	#10 counter$count = 72731;
	#10 counter$count = 72732;
	#10 counter$count = 72733;
	#10 counter$count = 72734;
	#10 counter$count = 72735;
	#10 counter$count = 72736;
	#10 counter$count = 72737;
	#10 counter$count = 72738;
	#10 counter$count = 72739;
	#10 counter$count = 72740;
	#10 counter$count = 72741;
	#10 counter$count = 72742;
	#10 counter$count = 72743;
	#10 counter$count = 72744;
	#10 counter$count = 72745;
	#10 counter$count = 72746;
	#10 counter$count = 72747;
	#10 counter$count = 72748;
	#10 counter$count = 72749;
	#10 counter$count = 72750;
	#10 counter$count = 72751;
	#10 counter$count = 72752;
	#10 counter$count = 72753;
	#10 counter$count = 72754;
	#10 counter$count = 72755;
	#10 counter$count = 72756;
	#10 counter$count = 72757;
	#10 counter$count = 72758;
	#10 counter$count = 72759;
	#10 counter$count = 72760;
	#10 counter$count = 72761;
	#10 counter$count = 72762;
	#10 counter$count = 72763;
	#10 counter$count = 72764;
	#10 counter$count = 72765;
	#10 counter$count = 72766;
	#10 counter$count = 72767;
	#10 counter$count = 72768;
	#10 counter$count = 72769;
	#10 counter$count = 72770;
	#10 counter$count = 72771;
	#10 counter$count = 72772;
	#10 counter$count = 72773;
	#10 counter$count = 72774;
	#10 counter$count = 72775;
	#10 counter$count = 72776;
	#10 counter$count = 72777;
	#10 counter$count = 72778;
	#10 counter$count = 72779;
	#10 counter$count = 72780;
	#10 counter$count = 72781;
	#10 counter$count = 72782;
	#10 counter$count = 72783;
	#10 counter$count = 72784;
	#10 counter$count = 72785;
	#10 counter$count = 72786;
	#10 counter$count = 72787;
	#10 counter$count = 72788;
	#10 counter$count = 72789;
	#10 counter$count = 72790;
	#10 counter$count = 72791;
	#10 counter$count = 72792;
	#10 counter$count = 72793;
	#10 counter$count = 72794;
	#10 counter$count = 72795;
	#10 counter$count = 72796;
	#10 counter$count = 72797;
	#10 counter$count = 72798;
	#10 counter$count = 72799;
	#10 counter$count = 72800;
	#10 counter$count = 72801;
	#10 counter$count = 72802;
	#10 counter$count = 72803;
	#10 counter$count = 72804;
	#10 counter$count = 72805;
	#10 counter$count = 72806;
	#10 counter$count = 72807;
	#10 counter$count = 72808;
	#10 counter$count = 72809;
	#10 counter$count = 72810;
	#10 counter$count = 72811;
	#10 counter$count = 72812;
	#10 counter$count = 72813;
	#10 counter$count = 72814;
	#10 counter$count = 72815;
	#10 counter$count = 72816;
	#10 counter$count = 72817;
	#10 counter$count = 72818;
	#10 counter$count = 72819;
	#10 counter$count = 72820;
	#10 counter$count = 72821;
	#10 counter$count = 72822;
	#10 counter$count = 72823;
	#10 counter$count = 72824;
	#10 counter$count = 72825;
	#10 counter$count = 72826;
	#10 counter$count = 72827;
	#10 counter$count = 72828;
	#10 counter$count = 72829;
	#10 counter$count = 72830;
	#10 counter$count = 72831;
	#10 counter$count = 72832;
	#10 counter$count = 72833;
	#10 counter$count = 72834;
	#10 counter$count = 72835;
	#10 counter$count = 72836;
	#10 counter$count = 72837;
	#10 counter$count = 72838;
	#10 counter$count = 72839;
	#10 counter$count = 72840;
	#10 counter$count = 72841;
	#10 counter$count = 72842;
	#10 counter$count = 72843;
	#10 counter$count = 72844;
	#10 counter$count = 72845;
	#10 counter$count = 72846;
	#10 counter$count = 72847;
	#10 counter$count = 72848;
	#10 counter$count = 72849;
	#10 counter$count = 72850;
	#10 counter$count = 72851;
	#10 counter$count = 72852;
	#10 counter$count = 72853;
	#10 counter$count = 72854;
	#10 counter$count = 72855;
	#10 counter$count = 72856;
	#10 counter$count = 72857;
	#10 counter$count = 72858;
	#10 counter$count = 72859;
	#10 counter$count = 72860;
	#10 counter$count = 72861;
	#10 counter$count = 72862;
	#10 counter$count = 72863;
	#10 counter$count = 72864;
	#10 counter$count = 72865;
	#10 counter$count = 72866;
	#10 counter$count = 72867;
	#10 counter$count = 72868;
	#10 counter$count = 72869;
	#10 counter$count = 72870;
	#10 counter$count = 72871;
	#10 counter$count = 72872;
	#10 counter$count = 72873;
	#10 counter$count = 72874;
	#10 counter$count = 72875;
	#10 counter$count = 72876;
	#10 counter$count = 72877;
	#10 counter$count = 72878;
	#10 counter$count = 72879;
	#10 counter$count = 72880;
	#10 counter$count = 72881;
	#10 counter$count = 72882;
	#10 counter$count = 72883;
	#10 counter$count = 72884;
	#10 counter$count = 72885;
	#10 counter$count = 72886;
	#10 counter$count = 72887;
	#10 counter$count = 72888;
	#10 counter$count = 72889;
	#10 counter$count = 72890;
	#10 counter$count = 72891;
	#10 counter$count = 72892;
	#10 counter$count = 72893;
	#10 counter$count = 72894;
	#10 counter$count = 72895;
	#10 counter$count = 72896;
	#10 counter$count = 72897;
	#10 counter$count = 72898;
	#10 counter$count = 72899;
	#10 counter$count = 72900;
	#10 counter$count = 72901;
	#10 counter$count = 72902;
	#10 counter$count = 72903;
	#10 counter$count = 72904;
	#10 counter$count = 72905;
	#10 counter$count = 72906;
	#10 counter$count = 72907;
	#10 counter$count = 72908;
	#10 counter$count = 72909;
	#10 counter$count = 72910;
	#10 counter$count = 72911;
	#10 counter$count = 72912;
	#10 counter$count = 72913;
	#10 counter$count = 72914;
	#10 counter$count = 72915;
	#10 counter$count = 72916;
	#10 counter$count = 72917;
	#10 counter$count = 72918;
	#10 counter$count = 72919;
	#10 counter$count = 72920;
	#10 counter$count = 72921;
	#10 counter$count = 72922;
	#10 counter$count = 72923;
	#10 counter$count = 72924;
	#10 counter$count = 72925;
	#10 counter$count = 72926;
	#10 counter$count = 72927;
	#10 counter$count = 72928;
	#10 counter$count = 72929;
	#10 counter$count = 72930;
	#10 counter$count = 72931;
	#10 counter$count = 72932;
	#10 counter$count = 72933;
	#10 counter$count = 72934;
	#10 counter$count = 72935;
	#10 counter$count = 72936;
	#10 counter$count = 72937;
	#10 counter$count = 72938;
	#10 counter$count = 72939;
	#10 counter$count = 72940;
	#10 counter$count = 72941;
	#10 counter$count = 72942;
	#10 counter$count = 72943;
	#10 counter$count = 72944;
	#10 counter$count = 72945;
	#10 counter$count = 72946;
	#10 counter$count = 72947;
	#10 counter$count = 72948;
	#10 counter$count = 72949;
	#10 counter$count = 72950;
	#10 counter$count = 72951;
	#10 counter$count = 72952;
	#10 counter$count = 72953;
	#10 counter$count = 72954;
	#10 counter$count = 72955;
	#10 counter$count = 72956;
	#10 counter$count = 72957;
	#10 counter$count = 72958;
	#10 counter$count = 72959;
	#10 counter$count = 72960;
	#10 counter$count = 72961;
	#10 counter$count = 72962;
	#10 counter$count = 72963;
	#10 counter$count = 72964;
	#10 counter$count = 72965;
	#10 counter$count = 72966;
	#10 counter$count = 72967;
	#10 counter$count = 72968;
	#10 counter$count = 72969;
	#10 counter$count = 72970;
	#10 counter$count = 72971;
	#10 counter$count = 72972;
	#10 counter$count = 72973;
	#10 counter$count = 72974;
	#10 counter$count = 72975;
	#10 counter$count = 72976;
	#10 counter$count = 72977;
	#10 counter$count = 72978;
	#10 counter$count = 72979;
	#10 counter$count = 72980;
	#10 counter$count = 72981;
	#10 counter$count = 72982;
	#10 counter$count = 72983;
	#10 counter$count = 72984;
	#10 counter$count = 72985;
	#10 counter$count = 72986;
	#10 counter$count = 72987;
	#10 counter$count = 72988;
	#10 counter$count = 72989;
	#10 counter$count = 72990;
	#10 counter$count = 72991;
	#10 counter$count = 72992;
	#10 counter$count = 72993;
	#10 counter$count = 72994;
	#10 counter$count = 72995;
	#10 counter$count = 72996;
	#10 counter$count = 72997;
	#10 counter$count = 72998;
	#10 counter$count = 72999;
	#10 counter$count = 73000;
	#10 counter$count = 73001;
	#10 counter$count = 73002;
	#10 counter$count = 73003;
	#10 counter$count = 73004;
	#10 counter$count = 73005;
	#10 counter$count = 73006;
	#10 counter$count = 73007;
	#10 counter$count = 73008;
	#10 counter$count = 73009;
	#10 counter$count = 73010;
	#10 counter$count = 73011;
	#10 counter$count = 73012;
	#10 counter$count = 73013;
	#10 counter$count = 73014;
	#10 counter$count = 73015;
	#10 counter$count = 73016;
	#10 counter$count = 73017;
	#10 counter$count = 73018;
	#10 counter$count = 73019;
	#10 counter$count = 73020;
	#10 counter$count = 73021;
	#10 counter$count = 73022;
	#10 counter$count = 73023;
	#10 counter$count = 73024;
	#10 counter$count = 73025;
	#10 counter$count = 73026;
	#10 counter$count = 73027;
	#10 counter$count = 73028;
	#10 counter$count = 73029;
	#10 counter$count = 73030;
	#10 counter$count = 73031;
	#10 counter$count = 73032;
	#10 counter$count = 73033;
	#10 counter$count = 73034;
	#10 counter$count = 73035;
	#10 counter$count = 73036;
	#10 counter$count = 73037;
	#10 counter$count = 73038;
	#10 counter$count = 73039;
	#10 counter$count = 73040;
	#10 counter$count = 73041;
	#10 counter$count = 73042;
	#10 counter$count = 73043;
	#10 counter$count = 73044;
	#10 counter$count = 73045;
	#10 counter$count = 73046;
	#10 counter$count = 73047;
	#10 counter$count = 73048;
	#10 counter$count = 73049;
	#10 counter$count = 73050;
	#10 counter$count = 73051;
	#10 counter$count = 73052;
	#10 counter$count = 73053;
	#10 counter$count = 73054;
	#10 counter$count = 73055;
	#10 counter$count = 73056;
	#10 counter$count = 73057;
	#10 counter$count = 73058;
	#10 counter$count = 73059;
	#10 counter$count = 73060;
	#10 counter$count = 73061;
	#10 counter$count = 73062;
	#10 counter$count = 73063;
	#10 counter$count = 73064;
	#10 counter$count = 73065;
	#10 counter$count = 73066;
	#10 counter$count = 73067;
	#10 counter$count = 73068;
	#10 counter$count = 73069;
	#10 counter$count = 73070;
	#10 counter$count = 73071;
	#10 counter$count = 73072;
	#10 counter$count = 73073;
	#10 counter$count = 73074;
	#10 counter$count = 73075;
	#10 counter$count = 73076;
	#10 counter$count = 73077;
	#10 counter$count = 73078;
	#10 counter$count = 73079;
	#10 counter$count = 73080;
	#10 counter$count = 73081;
	#10 counter$count = 73082;
	#10 counter$count = 73083;
	#10 counter$count = 73084;
	#10 counter$count = 73085;
	#10 counter$count = 73086;
	#10 counter$count = 73087;
	#10 counter$count = 73088;
	#10 counter$count = 73089;
	#10 counter$count = 73090;
	#10 counter$count = 73091;
	#10 counter$count = 73092;
	#10 counter$count = 73093;
	#10 counter$count = 73094;
	#10 counter$count = 73095;
	#10 counter$count = 73096;
	#10 counter$count = 73097;
	#10 counter$count = 73098;
	#10 counter$count = 73099;
	#10 counter$count = 73100;
	#10 counter$count = 73101;
	#10 counter$count = 73102;
	#10 counter$count = 73103;
	#10 counter$count = 73104;
	#10 counter$count = 73105;
	#10 counter$count = 73106;
	#10 counter$count = 73107;
	#10 counter$count = 73108;
	#10 counter$count = 73109;
	#10 counter$count = 73110;
	#10 counter$count = 73111;
	#10 counter$count = 73112;
	#10 counter$count = 73113;
	#10 counter$count = 73114;
	#10 counter$count = 73115;
	#10 counter$count = 73116;
	#10 counter$count = 73117;
	#10 counter$count = 73118;
	#10 counter$count = 73119;
	#10 counter$count = 73120;
	#10 counter$count = 73121;
	#10 counter$count = 73122;
	#10 counter$count = 73123;
	#10 counter$count = 73124;
	#10 counter$count = 73125;
	#10 counter$count = 73126;
	#10 counter$count = 73127;
	#10 counter$count = 73128;
	#10 counter$count = 73129;
	#10 counter$count = 73130;
	#10 counter$count = 73131;
	#10 counter$count = 73132;
	#10 counter$count = 73133;
	#10 counter$count = 73134;
	#10 counter$count = 73135;
	#10 counter$count = 73136;
	#10 counter$count = 73137;
	#10 counter$count = 73138;
	#10 counter$count = 73139;
	#10 counter$count = 73140;
	#10 counter$count = 73141;
	#10 counter$count = 73142;
	#10 counter$count = 73143;
	#10 counter$count = 73144;
	#10 counter$count = 73145;
	#10 counter$count = 73146;
	#10 counter$count = 73147;
	#10 counter$count = 73148;
	#10 counter$count = 73149;
	#10 counter$count = 73150;
	#10 counter$count = 73151;
	#10 counter$count = 73152;
	#10 counter$count = 73153;
	#10 counter$count = 73154;
	#10 counter$count = 73155;
	#10 counter$count = 73156;
	#10 counter$count = 73157;
	#10 counter$count = 73158;
	#10 counter$count = 73159;
	#10 counter$count = 73160;
	#10 counter$count = 73161;
	#10 counter$count = 73162;
	#10 counter$count = 73163;
	#10 counter$count = 73164;
	#10 counter$count = 73165;
	#10 counter$count = 73166;
	#10 counter$count = 73167;
	#10 counter$count = 73168;
	#10 counter$count = 73169;
	#10 counter$count = 73170;
	#10 counter$count = 73171;
	#10 counter$count = 73172;
	#10 counter$count = 73173;
	#10 counter$count = 73174;
	#10 counter$count = 73175;
	#10 counter$count = 73176;
	#10 counter$count = 73177;
	#10 counter$count = 73178;
	#10 counter$count = 73179;
	#10 counter$count = 73180;
	#10 counter$count = 73181;
	#10 counter$count = 73182;
	#10 counter$count = 73183;
	#10 counter$count = 73184;
	#10 counter$count = 73185;
	#10 counter$count = 73186;
	#10 counter$count = 73187;
	#10 counter$count = 73188;
	#10 counter$count = 73189;
	#10 counter$count = 73190;
	#10 counter$count = 73191;
	#10 counter$count = 73192;
	#10 counter$count = 73193;
	#10 counter$count = 73194;
	#10 counter$count = 73195;
	#10 counter$count = 73196;
	#10 counter$count = 73197;
	#10 counter$count = 73198;
	#10 counter$count = 73199;
	#10 counter$count = 73200;
	#10 counter$count = 73201;
	#10 counter$count = 73202;
	#10 counter$count = 73203;
	#10 counter$count = 73204;
	#10 counter$count = 73205;
	#10 counter$count = 73206;
	#10 counter$count = 73207;
	#10 counter$count = 73208;
	#10 counter$count = 73209;
	#10 counter$count = 73210;
	#10 counter$count = 73211;
	#10 counter$count = 73212;
	#10 counter$count = 73213;
	#10 counter$count = 73214;
	#10 counter$count = 73215;
	#10 counter$count = 73216;
	#10 counter$count = 73217;
	#10 counter$count = 73218;
	#10 counter$count = 73219;
	#10 counter$count = 73220;
	#10 counter$count = 73221;
	#10 counter$count = 73222;
	#10 counter$count = 73223;
	#10 counter$count = 73224;
	#10 counter$count = 73225;
	#10 counter$count = 73226;
	#10 counter$count = 73227;
	#10 counter$count = 73228;
	#10 counter$count = 73229;
	#10 counter$count = 73230;
	#10 counter$count = 73231;
	#10 counter$count = 73232;
	#10 counter$count = 73233;
	#10 counter$count = 73234;
	#10 counter$count = 73235;
	#10 counter$count = 73236;
	#10 counter$count = 73237;
	#10 counter$count = 73238;
	#10 counter$count = 73239;
	#10 counter$count = 73240;
	#10 counter$count = 73241;
	#10 counter$count = 73242;
	#10 counter$count = 73243;
	#10 counter$count = 73244;
	#10 counter$count = 73245;
	#10 counter$count = 73246;
	#10 counter$count = 73247;
	#10 counter$count = 73248;
	#10 counter$count = 73249;
	#10 counter$count = 73250;
	#10 counter$count = 73251;
	#10 counter$count = 73252;
	#10 counter$count = 73253;
	#10 counter$count = 73254;
	#10 counter$count = 73255;
	#10 counter$count = 73256;
	#10 counter$count = 73257;
	#10 counter$count = 73258;
	#10 counter$count = 73259;
	#10 counter$count = 73260;
	#10 counter$count = 73261;
	#10 counter$count = 73262;
	#10 counter$count = 73263;
	#10 counter$count = 73264;
	#10 counter$count = 73265;
	#10 counter$count = 73266;
	#10 counter$count = 73267;
	#10 counter$count = 73268;
	#10 counter$count = 73269;
	#10 counter$count = 73270;
	#10 counter$count = 73271;
	#10 counter$count = 73272;
	#10 counter$count = 73273;
	#10 counter$count = 73274;
	#10 counter$count = 73275;
	#10 counter$count = 73276;
	#10 counter$count = 73277;
	#10 counter$count = 73278;
	#10 counter$count = 73279;
	#10 counter$count = 73280;
	#10 counter$count = 73281;
	#10 counter$count = 73282;
	#10 counter$count = 73283;
	#10 counter$count = 73284;
	#10 counter$count = 73285;
	#10 counter$count = 73286;
	#10 counter$count = 73287;
	#10 counter$count = 73288;
	#10 counter$count = 73289;
	#10 counter$count = 73290;
	#10 counter$count = 73291;
	#10 counter$count = 73292;
	#10 counter$count = 73293;
	#10 counter$count = 73294;
	#10 counter$count = 73295;
	#10 counter$count = 73296;
	#10 counter$count = 73297;
	#10 counter$count = 73298;
	#10 counter$count = 73299;
	#10 counter$count = 73300;
	#10 counter$count = 73301;
	#10 counter$count = 73302;
	#10 counter$count = 73303;
	#10 counter$count = 73304;
	#10 counter$count = 73305;
	#10 counter$count = 73306;
	#10 counter$count = 73307;
	#10 counter$count = 73308;
	#10 counter$count = 73309;
	#10 counter$count = 73310;
	#10 counter$count = 73311;
	#10 counter$count = 73312;
	#10 counter$count = 73313;
	#10 counter$count = 73314;
	#10 counter$count = 73315;
	#10 counter$count = 73316;
	#10 counter$count = 73317;
	#10 counter$count = 73318;
	#10 counter$count = 73319;
	#10 counter$count = 73320;
	#10 counter$count = 73321;
	#10 counter$count = 73322;
	#10 counter$count = 73323;
	#10 counter$count = 73324;
	#10 counter$count = 73325;
	#10 counter$count = 73326;
	#10 counter$count = 73327;
	#10 counter$count = 73328;
	#10 counter$count = 73329;
	#10 counter$count = 73330;
	#10 counter$count = 73331;
	#10 counter$count = 73332;
	#10 counter$count = 73333;
	#10 counter$count = 73334;
	#10 counter$count = 73335;
	#10 counter$count = 73336;
	#10 counter$count = 73337;
	#10 counter$count = 73338;
	#10 counter$count = 73339;
	#10 counter$count = 73340;
	#10 counter$count = 73341;
	#10 counter$count = 73342;
	#10 counter$count = 73343;
	#10 counter$count = 73344;
	#10 counter$count = 73345;
	#10 counter$count = 73346;
	#10 counter$count = 73347;
	#10 counter$count = 73348;
	#10 counter$count = 73349;
	#10 counter$count = 73350;
	#10 counter$count = 73351;
	#10 counter$count = 73352;
	#10 counter$count = 73353;
	#10 counter$count = 73354;
	#10 counter$count = 73355;
	#10 counter$count = 73356;
	#10 counter$count = 73357;
	#10 counter$count = 73358;
	#10 counter$count = 73359;
	#10 counter$count = 73360;
	#10 counter$count = 73361;
	#10 counter$count = 73362;
	#10 counter$count = 73363;
	#10 counter$count = 73364;
	#10 counter$count = 73365;
	#10 counter$count = 73366;
	#10 counter$count = 73367;
	#10 counter$count = 73368;
	#10 counter$count = 73369;
	#10 counter$count = 73370;
	#10 counter$count = 73371;
	#10 counter$count = 73372;
	#10 counter$count = 73373;
	#10 counter$count = 73374;
	#10 counter$count = 73375;
	#10 counter$count = 73376;
	#10 counter$count = 73377;
	#10 counter$count = 73378;
	#10 counter$count = 73379;
	#10 counter$count = 73380;
	#10 counter$count = 73381;
	#10 counter$count = 73382;
	#10 counter$count = 73383;
	#10 counter$count = 73384;
	#10 counter$count = 73385;
	#10 counter$count = 73386;
	#10 counter$count = 73387;
	#10 counter$count = 73388;
	#10 counter$count = 73389;
	#10 counter$count = 73390;
	#10 counter$count = 73391;
	#10 counter$count = 73392;
	#10 counter$count = 73393;
	#10 counter$count = 73394;
	#10 counter$count = 73395;
	#10 counter$count = 73396;
	#10 counter$count = 73397;
	#10 counter$count = 73398;
	#10 counter$count = 73399;
	#10 counter$count = 73400;
	#10 counter$count = 73401;
	#10 counter$count = 73402;
	#10 counter$count = 73403;
	#10 counter$count = 73404;
	#10 counter$count = 73405;
	#10 counter$count = 73406;
	#10 counter$count = 73407;
	#10 counter$count = 73408;
	#10 counter$count = 73409;
	#10 counter$count = 73410;
	#10 counter$count = 73411;
	#10 counter$count = 73412;
	#10 counter$count = 73413;
	#10 counter$count = 73414;
	#10 counter$count = 73415;
	#10 counter$count = 73416;
	#10 counter$count = 73417;
	#10 counter$count = 73418;
	#10 counter$count = 73419;
	#10 counter$count = 73420;
	#10 counter$count = 73421;
	#10 counter$count = 73422;
	#10 counter$count = 73423;
	#10 counter$count = 73424;
	#10 counter$count = 73425;
	#10 counter$count = 73426;
	#10 counter$count = 73427;
	#10 counter$count = 73428;
	#10 counter$count = 73429;
	#10 counter$count = 73430;
	#10 counter$count = 73431;
	#10 counter$count = 73432;
	#10 counter$count = 73433;
	#10 counter$count = 73434;
	#10 counter$count = 73435;
	#10 counter$count = 73436;
	#10 counter$count = 73437;
	#10 counter$count = 73438;
	#10 counter$count = 73439;
	#10 counter$count = 73440;
	#10 counter$count = 73441;
	#10 counter$count = 73442;
	#10 counter$count = 73443;
	#10 counter$count = 73444;
	#10 counter$count = 73445;
	#10 counter$count = 73446;
	#10 counter$count = 73447;
	#10 counter$count = 73448;
	#10 counter$count = 73449;
	#10 counter$count = 73450;
	#10 counter$count = 73451;
	#10 counter$count = 73452;
	#10 counter$count = 73453;
	#10 counter$count = 73454;
	#10 counter$count = 73455;
	#10 counter$count = 73456;
	#10 counter$count = 73457;
	#10 counter$count = 73458;
	#10 counter$count = 73459;
	#10 counter$count = 73460;
	#10 counter$count = 73461;
	#10 counter$count = 73462;
	#10 counter$count = 73463;
	#10 counter$count = 73464;
	#10 counter$count = 73465;
	#10 counter$count = 73466;
	#10 counter$count = 73467;
	#10 counter$count = 73468;
	#10 counter$count = 73469;
	#10 counter$count = 73470;
	#10 counter$count = 73471;
	#10 counter$count = 73472;
	#10 counter$count = 73473;
	#10 counter$count = 73474;
	#10 counter$count = 73475;
	#10 counter$count = 73476;
	#10 counter$count = 73477;
	#10 counter$count = 73478;
	#10 counter$count = 73479;
	#10 counter$count = 73480;
	#10 counter$count = 73481;
	#10 counter$count = 73482;
	#10 counter$count = 73483;
	#10 counter$count = 73484;
	#10 counter$count = 73485;
	#10 counter$count = 73486;
	#10 counter$count = 73487;
	#10 counter$count = 73488;
	#10 counter$count = 73489;
	#10 counter$count = 73490;
	#10 counter$count = 73491;
	#10 counter$count = 73492;
	#10 counter$count = 73493;
	#10 counter$count = 73494;
	#10 counter$count = 73495;
	#10 counter$count = 73496;
	#10 counter$count = 73497;
	#10 counter$count = 73498;
	#10 counter$count = 73499;
	#10 counter$count = 73500;
	#10 counter$count = 73501;
	#10 counter$count = 73502;
	#10 counter$count = 73503;
	#10 counter$count = 73504;
	#10 counter$count = 73505;
	#10 counter$count = 73506;
	#10 counter$count = 73507;
	#10 counter$count = 73508;
	#10 counter$count = 73509;
	#10 counter$count = 73510;
	#10 counter$count = 73511;
	#10 counter$count = 73512;
	#10 counter$count = 73513;
	#10 counter$count = 73514;
	#10 counter$count = 73515;
	#10 counter$count = 73516;
	#10 counter$count = 73517;
	#10 counter$count = 73518;
	#10 counter$count = 73519;
	#10 counter$count = 73520;
	#10 counter$count = 73521;
	#10 counter$count = 73522;
	#10 counter$count = 73523;
	#10 counter$count = 73524;
	#10 counter$count = 73525;
	#10 counter$count = 73526;
	#10 counter$count = 73527;
	#10 counter$count = 73528;
	#10 counter$count = 73529;
	#10 counter$count = 73530;
	#10 counter$count = 73531;
	#10 counter$count = 73532;
	#10 counter$count = 73533;
	#10 counter$count = 73534;
	#10 counter$count = 73535;
	#10 counter$count = 73536;
	#10 counter$count = 73537;
	#10 counter$count = 73538;
	#10 counter$count = 73539;
	#10 counter$count = 73540;
	#10 counter$count = 73541;
	#10 counter$count = 73542;
	#10 counter$count = 73543;
	#10 counter$count = 73544;
	#10 counter$count = 73545;
	#10 counter$count = 73546;
	#10 counter$count = 73547;
	#10 counter$count = 73548;
	#10 counter$count = 73549;
	#10 counter$count = 73550;
	#10 counter$count = 73551;
	#10 counter$count = 73552;
	#10 counter$count = 73553;
	#10 counter$count = 73554;
	#10 counter$count = 73555;
	#10 counter$count = 73556;
	#10 counter$count = 73557;
	#10 counter$count = 73558;
	#10 counter$count = 73559;
	#10 counter$count = 73560;
	#10 counter$count = 73561;
	#10 counter$count = 73562;
	#10 counter$count = 73563;
	#10 counter$count = 73564;
	#10 counter$count = 73565;
	#10 counter$count = 73566;
	#10 counter$count = 73567;
	#10 counter$count = 73568;
	#10 counter$count = 73569;
	#10 counter$count = 73570;
	#10 counter$count = 73571;
	#10 counter$count = 73572;
	#10 counter$count = 73573;
	#10 counter$count = 73574;
	#10 counter$count = 73575;
	#10 counter$count = 73576;
	#10 counter$count = 73577;
	#10 counter$count = 73578;
	#10 counter$count = 73579;
	#10 counter$count = 73580;
	#10 counter$count = 73581;
	#10 counter$count = 73582;
	#10 counter$count = 73583;
	#10 counter$count = 73584;
	#10 counter$count = 73585;
	#10 counter$count = 73586;
	#10 counter$count = 73587;
	#10 counter$count = 73588;
	#10 counter$count = 73589;
	#10 counter$count = 73590;
	#10 counter$count = 73591;
	#10 counter$count = 73592;
	#10 counter$count = 73593;
	#10 counter$count = 73594;
	#10 counter$count = 73595;
	#10 counter$count = 73596;
	#10 counter$count = 73597;
	#10 counter$count = 73598;
	#10 counter$count = 73599;
	#10 counter$count = 73600;
	#10 counter$count = 73601;
	#10 counter$count = 73602;
	#10 counter$count = 73603;
	#10 counter$count = 73604;
	#10 counter$count = 73605;
	#10 counter$count = 73606;
	#10 counter$count = 73607;
	#10 counter$count = 73608;
	#10 counter$count = 73609;
	#10 counter$count = 73610;
	#10 counter$count = 73611;
	#10 counter$count = 73612;
	#10 counter$count = 73613;
	#10 counter$count = 73614;
	#10 counter$count = 73615;
	#10 counter$count = 73616;
	#10 counter$count = 73617;
	#10 counter$count = 73618;
	#10 counter$count = 73619;
	#10 counter$count = 73620;
	#10 counter$count = 73621;
	#10 counter$count = 73622;
	#10 counter$count = 73623;
	#10 counter$count = 73624;
	#10 counter$count = 73625;
	#10 counter$count = 73626;
	#10 counter$count = 73627;
	#10 counter$count = 73628;
	#10 counter$count = 73629;
	#10 counter$count = 73630;
	#10 counter$count = 73631;
	#10 counter$count = 73632;
	#10 counter$count = 73633;
	#10 counter$count = 73634;
	#10 counter$count = 73635;
	#10 counter$count = 73636;
	#10 counter$count = 73637;
	#10 counter$count = 73638;
	#10 counter$count = 73639;
	#10 counter$count = 73640;
	#10 counter$count = 73641;
	#10 counter$count = 73642;
	#10 counter$count = 73643;
	#10 counter$count = 73644;
	#10 counter$count = 73645;
	#10 counter$count = 73646;
	#10 counter$count = 73647;
	#10 counter$count = 73648;
	#10 counter$count = 73649;
	#10 counter$count = 73650;
	#10 counter$count = 73651;
	#10 counter$count = 73652;
	#10 counter$count = 73653;
	#10 counter$count = 73654;
	#10 counter$count = 73655;
	#10 counter$count = 73656;
	#10 counter$count = 73657;
	#10 counter$count = 73658;
	#10 counter$count = 73659;
	#10 counter$count = 73660;
	#10 counter$count = 73661;
	#10 counter$count = 73662;
	#10 counter$count = 73663;
	#10 counter$count = 73664;
	#10 counter$count = 73665;
	#10 counter$count = 73666;
	#10 counter$count = 73667;
	#10 counter$count = 73668;
	#10 counter$count = 73669;
	#10 counter$count = 73670;
	#10 counter$count = 73671;
	#10 counter$count = 73672;
	#10 counter$count = 73673;
	#10 counter$count = 73674;
	#10 counter$count = 73675;
	#10 counter$count = 73676;
	#10 counter$count = 73677;
	#10 counter$count = 73678;
	#10 counter$count = 73679;
	#10 counter$count = 73680;
	#10 counter$count = 73681;
	#10 counter$count = 73682;
	#10 counter$count = 73683;
	#10 counter$count = 73684;
	#10 counter$count = 73685;
	#10 counter$count = 73686;
	#10 counter$count = 73687;
	#10 counter$count = 73688;
	#10 counter$count = 73689;
	#10 counter$count = 73690;
	#10 counter$count = 73691;
	#10 counter$count = 73692;
	#10 counter$count = 73693;
	#10 counter$count = 73694;
	#10 counter$count = 73695;
	#10 counter$count = 73696;
	#10 counter$count = 73697;
	#10 counter$count = 73698;
	#10 counter$count = 73699;
	#10 counter$count = 73700;
	#10 counter$count = 73701;
	#10 counter$count = 73702;
	#10 counter$count = 73703;
	#10 counter$count = 73704;
	#10 counter$count = 73705;
	#10 counter$count = 73706;
	#10 counter$count = 73707;
	#10 counter$count = 73708;
	#10 counter$count = 73709;
	#10 counter$count = 73710;
	#10 counter$count = 73711;
	#10 counter$count = 73712;
	#10 counter$count = 73713;
	#10 counter$count = 73714;
	#10 counter$count = 73715;
	#10 counter$count = 73716;
	#10 counter$count = 73717;
	#10 counter$count = 73718;
	#10 counter$count = 73719;
	#10 counter$count = 73720;
	#10 counter$count = 73721;
	#10 counter$count = 73722;
	#10 counter$count = 73723;
	#10 counter$count = 73724;
	#10 counter$count = 73725;
	#10 counter$count = 73726;
	#10 counter$count = 73727;
	#10 counter$count = 73728;
	#10 counter$count = 73729;
	#10 counter$count = 73730;
	#10 counter$count = 73731;
	#10 counter$count = 73732;
	#10 counter$count = 73733;
	#10 counter$count = 73734;
	#10 counter$count = 73735;
	#10 counter$count = 73736;
	#10 counter$count = 73737;
	#10 counter$count = 73738;
	#10 counter$count = 73739;
	#10 counter$count = 73740;
	#10 counter$count = 73741;
	#10 counter$count = 73742;
	#10 counter$count = 73743;
	#10 counter$count = 73744;
	#10 counter$count = 73745;
	#10 counter$count = 73746;
	#10 counter$count = 73747;
	#10 counter$count = 73748;
	#10 counter$count = 73749;
	#10 counter$count = 73750;
	#10 counter$count = 73751;
	#10 counter$count = 73752;
	#10 counter$count = 73753;
	#10 counter$count = 73754;
	#10 counter$count = 73755;
	#10 counter$count = 73756;
	#10 counter$count = 73757;
	#10 counter$count = 73758;
	#10 counter$count = 73759;
	#10 counter$count = 73760;
	#10 counter$count = 73761;
	#10 counter$count = 73762;
	#10 counter$count = 73763;
	#10 counter$count = 73764;
	#10 counter$count = 73765;
	#10 counter$count = 73766;
	#10 counter$count = 73767;
	#10 counter$count = 73768;
	#10 counter$count = 73769;
	#10 counter$count = 73770;
	#10 counter$count = 73771;
	#10 counter$count = 73772;
	#10 counter$count = 73773;
	#10 counter$count = 73774;
	#10 counter$count = 73775;
	#10 counter$count = 73776;
	#10 counter$count = 73777;
	#10 counter$count = 73778;
	#10 counter$count = 73779;
	#10 counter$count = 73780;
	#10 counter$count = 73781;
	#10 counter$count = 73782;
	#10 counter$count = 73783;
	#10 counter$count = 73784;
	#10 counter$count = 73785;
	#10 counter$count = 73786;
	#10 counter$count = 73787;
	#10 counter$count = 73788;
	#10 counter$count = 73789;
	#10 counter$count = 73790;
	#10 counter$count = 73791;
	#10 counter$count = 73792;
	#10 counter$count = 73793;
	#10 counter$count = 73794;
	#10 counter$count = 73795;
	#10 counter$count = 73796;
	#10 counter$count = 73797;
	#10 counter$count = 73798;
	#10 counter$count = 73799;
	#10 counter$count = 73800;
	#10 counter$count = 73801;
	#10 counter$count = 73802;
	#10 counter$count = 73803;
	#10 counter$count = 73804;
	#10 counter$count = 73805;
	#10 counter$count = 73806;
	#10 counter$count = 73807;
	#10 counter$count = 73808;
	#10 counter$count = 73809;
	#10 counter$count = 73810;
	#10 counter$count = 73811;
	#10 counter$count = 73812;
	#10 counter$count = 73813;
	#10 counter$count = 73814;
	#10 counter$count = 73815;
	#10 counter$count = 73816;
	#10 counter$count = 73817;
	#10 counter$count = 73818;
	#10 counter$count = 73819;
	#10 counter$count = 73820;
	#10 counter$count = 73821;
	#10 counter$count = 73822;
	#10 counter$count = 73823;
	#10 counter$count = 73824;
	#10 counter$count = 73825;
	#10 counter$count = 73826;
	#10 counter$count = 73827;
	#10 counter$count = 73828;
	#10 counter$count = 73829;
	#10 counter$count = 73830;
	#10 counter$count = 73831;
	#10 counter$count = 73832;
	#10 counter$count = 73833;
	#10 counter$count = 73834;
	#10 counter$count = 73835;
	#10 counter$count = 73836;
	#10 counter$count = 73837;
	#10 counter$count = 73838;
	#10 counter$count = 73839;
	#10 counter$count = 73840;
	#10 counter$count = 73841;
	#10 counter$count = 73842;
	#10 counter$count = 73843;
	#10 counter$count = 73844;
	#10 counter$count = 73845;
	#10 counter$count = 73846;
	#10 counter$count = 73847;
	#10 counter$count = 73848;
	#10 counter$count = 73849;
	#10 counter$count = 73850;
	#10 counter$count = 73851;
	#10 counter$count = 73852;
	#10 counter$count = 73853;
	#10 counter$count = 73854;
	#10 counter$count = 73855;
	#10 counter$count = 73856;
	#10 counter$count = 73857;
	#10 counter$count = 73858;
	#10 counter$count = 73859;
	#10 counter$count = 73860;
	#10 counter$count = 73861;
	#10 counter$count = 73862;
	#10 counter$count = 73863;
	#10 counter$count = 73864;
	#10 counter$count = 73865;
	#10 counter$count = 73866;
	#10 counter$count = 73867;
	#10 counter$count = 73868;
	#10 counter$count = 73869;
	#10 counter$count = 73870;
	#10 counter$count = 73871;
	#10 counter$count = 73872;
	#10 counter$count = 73873;
	#10 counter$count = 73874;
	#10 counter$count = 73875;
	#10 counter$count = 73876;
	#10 counter$count = 73877;
	#10 counter$count = 73878;
	#10 counter$count = 73879;
	#10 counter$count = 73880;
	#10 counter$count = 73881;
	#10 counter$count = 73882;
	#10 counter$count = 73883;
	#10 counter$count = 73884;
	#10 counter$count = 73885;
	#10 counter$count = 73886;
	#10 counter$count = 73887;
	#10 counter$count = 73888;
	#10 counter$count = 73889;
	#10 counter$count = 73890;
	#10 counter$count = 73891;
	#10 counter$count = 73892;
	#10 counter$count = 73893;
	#10 counter$count = 73894;
	#10 counter$count = 73895;
	#10 counter$count = 73896;
	#10 counter$count = 73897;
	#10 counter$count = 73898;
	#10 counter$count = 73899;
	#10 counter$count = 73900;
	#10 counter$count = 73901;
	#10 counter$count = 73902;
	#10 counter$count = 73903;
	#10 counter$count = 73904;
	#10 counter$count = 73905;
	#10 counter$count = 73906;
	#10 counter$count = 73907;
	#10 counter$count = 73908;
	#10 counter$count = 73909;
	#10 counter$count = 73910;
	#10 counter$count = 73911;
	#10 counter$count = 73912;
	#10 counter$count = 73913;
	#10 counter$count = 73914;
	#10 counter$count = 73915;
	#10 counter$count = 73916;
	#10 counter$count = 73917;
	#10 counter$count = 73918;
	#10 counter$count = 73919;
	#10 counter$count = 73920;
	#10 counter$count = 73921;
	#10 counter$count = 73922;
	#10 counter$count = 73923;
	#10 counter$count = 73924;
	#10 counter$count = 73925;
	#10 counter$count = 73926;
	#10 counter$count = 73927;
	#10 counter$count = 73928;
	#10 counter$count = 73929;
	#10 counter$count = 73930;
	#10 counter$count = 73931;
	#10 counter$count = 73932;
	#10 counter$count = 73933;
	#10 counter$count = 73934;
	#10 counter$count = 73935;
	#10 counter$count = 73936;
	#10 counter$count = 73937;
	#10 counter$count = 73938;
	#10 counter$count = 73939;
	#10 counter$count = 73940;
	#10 counter$count = 73941;
	#10 counter$count = 73942;
	#10 counter$count = 73943;
	#10 counter$count = 73944;
	#10 counter$count = 73945;
	#10 counter$count = 73946;
	#10 counter$count = 73947;
	#10 counter$count = 73948;
	#10 counter$count = 73949;
	#10 counter$count = 73950;
	#10 counter$count = 73951;
	#10 counter$count = 73952;
	#10 counter$count = 73953;
	#10 counter$count = 73954;
	#10 counter$count = 73955;
	#10 counter$count = 73956;
	#10 counter$count = 73957;
	#10 counter$count = 73958;
	#10 counter$count = 73959;
	#10 counter$count = 73960;
	#10 counter$count = 73961;
	#10 counter$count = 73962;
	#10 counter$count = 73963;
	#10 counter$count = 73964;
	#10 counter$count = 73965;
	#10 counter$count = 73966;
	#10 counter$count = 73967;
	#10 counter$count = 73968;
	#10 counter$count = 73969;
	#10 counter$count = 73970;
	#10 counter$count = 73971;
	#10 counter$count = 73972;
	#10 counter$count = 73973;
	#10 counter$count = 73974;
	#10 counter$count = 73975;
	#10 counter$count = 73976;
	#10 counter$count = 73977;
	#10 counter$count = 73978;
	#10 counter$count = 73979;
	#10 counter$count = 73980;
	#10 counter$count = 73981;
	#10 counter$count = 73982;
	#10 counter$count = 73983;
	#10 counter$count = 73984;
	#10 counter$count = 73985;
	#10 counter$count = 73986;
	#10 counter$count = 73987;
	#10 counter$count = 73988;
	#10 counter$count = 73989;
	#10 counter$count = 73990;
	#10 counter$count = 73991;
	#10 counter$count = 73992;
	#10 counter$count = 73993;
	#10 counter$count = 73994;
	#10 counter$count = 73995;
	#10 counter$count = 73996;
	#10 counter$count = 73997;
	#10 counter$count = 73998;
	#10 counter$count = 73999;
	#10 counter$count = 74000;
	#10 counter$count = 74001;
	#10 counter$count = 74002;
	#10 counter$count = 74003;
	#10 counter$count = 74004;
	#10 counter$count = 74005;
	#10 counter$count = 74006;
	#10 counter$count = 74007;
	#10 counter$count = 74008;
	#10 counter$count = 74009;
	#10 counter$count = 74010;
	#10 counter$count = 74011;
	#10 counter$count = 74012;
	#10 counter$count = 74013;
	#10 counter$count = 74014;
	#10 counter$count = 74015;
	#10 counter$count = 74016;
	#10 counter$count = 74017;
	#10 counter$count = 74018;
	#10 counter$count = 74019;
	#10 counter$count = 74020;
	#10 counter$count = 74021;
	#10 counter$count = 74022;
	#10 counter$count = 74023;
	#10 counter$count = 74024;
	#10 counter$count = 74025;
	#10 counter$count = 74026;
	#10 counter$count = 74027;
	#10 counter$count = 74028;
	#10 counter$count = 74029;
	#10 counter$count = 74030;
	#10 counter$count = 74031;
	#10 counter$count = 74032;
	#10 counter$count = 74033;
	#10 counter$count = 74034;
	#10 counter$count = 74035;
	#10 counter$count = 74036;
	#10 counter$count = 74037;
	#10 counter$count = 74038;
	#10 counter$count = 74039;
	#10 counter$count = 74040;
	#10 counter$count = 74041;
	#10 counter$count = 74042;
	#10 counter$count = 74043;
	#10 counter$count = 74044;
	#10 counter$count = 74045;
	#10 counter$count = 74046;
	#10 counter$count = 74047;
	#10 counter$count = 74048;
	#10 counter$count = 74049;
	#10 counter$count = 74050;
	#10 counter$count = 74051;
	#10 counter$count = 74052;
	#10 counter$count = 74053;
	#10 counter$count = 74054;
	#10 counter$count = 74055;
	#10 counter$count = 74056;
	#10 counter$count = 74057;
	#10 counter$count = 74058;
	#10 counter$count = 74059;
	#10 counter$count = 74060;
	#10 counter$count = 74061;
	#10 counter$count = 74062;
	#10 counter$count = 74063;
	#10 counter$count = 74064;
	#10 counter$count = 74065;
	#10 counter$count = 74066;
	#10 counter$count = 74067;
	#10 counter$count = 74068;
	#10 counter$count = 74069;
	#10 counter$count = 74070;
	#10 counter$count = 74071;
	#10 counter$count = 74072;
	#10 counter$count = 74073;
	#10 counter$count = 74074;
	#10 counter$count = 74075;
	#10 counter$count = 74076;
	#10 counter$count = 74077;
	#10 counter$count = 74078;
	#10 counter$count = 74079;
	#10 counter$count = 74080;
	#10 counter$count = 74081;
	#10 counter$count = 74082;
	#10 counter$count = 74083;
	#10 counter$count = 74084;
	#10 counter$count = 74085;
	#10 counter$count = 74086;
	#10 counter$count = 74087;
	#10 counter$count = 74088;
	#10 counter$count = 74089;
	#10 counter$count = 74090;
	#10 counter$count = 74091;
	#10 counter$count = 74092;
	#10 counter$count = 74093;
	#10 counter$count = 74094;
	#10 counter$count = 74095;
	#10 counter$count = 74096;
	#10 counter$count = 74097;
	#10 counter$count = 74098;
	#10 counter$count = 74099;
	#10 counter$count = 74100;
	#10 counter$count = 74101;
	#10 counter$count = 74102;
	#10 counter$count = 74103;
	#10 counter$count = 74104;
	#10 counter$count = 74105;
	#10 counter$count = 74106;
	#10 counter$count = 74107;
	#10 counter$count = 74108;
	#10 counter$count = 74109;
	#10 counter$count = 74110;
	#10 counter$count = 74111;
	#10 counter$count = 74112;
	#10 counter$count = 74113;
	#10 counter$count = 74114;
	#10 counter$count = 74115;
	#10 counter$count = 74116;
	#10 counter$count = 74117;
	#10 counter$count = 74118;
	#10 counter$count = 74119;
	#10 counter$count = 74120;
	#10 counter$count = 74121;
	#10 counter$count = 74122;
	#10 counter$count = 74123;
	#10 counter$count = 74124;
	#10 counter$count = 74125;
	#10 counter$count = 74126;
	#10 counter$count = 74127;
	#10 counter$count = 74128;
	#10 counter$count = 74129;
	#10 counter$count = 74130;
	#10 counter$count = 74131;
	#10 counter$count = 74132;
	#10 counter$count = 74133;
	#10 counter$count = 74134;
	#10 counter$count = 74135;
	#10 counter$count = 74136;
	#10 counter$count = 74137;
	#10 counter$count = 74138;
	#10 counter$count = 74139;
	#10 counter$count = 74140;
	#10 counter$count = 74141;
	#10 counter$count = 74142;
	#10 counter$count = 74143;
	#10 counter$count = 74144;
	#10 counter$count = 74145;
	#10 counter$count = 74146;
	#10 counter$count = 74147;
	#10 counter$count = 74148;
	#10 counter$count = 74149;
	#10 counter$count = 74150;
	#10 counter$count = 74151;
	#10 counter$count = 74152;
	#10 counter$count = 74153;
	#10 counter$count = 74154;
	#10 counter$count = 74155;
	#10 counter$count = 74156;
	#10 counter$count = 74157;
	#10 counter$count = 74158;
	#10 counter$count = 74159;
	#10 counter$count = 74160;
	#10 counter$count = 74161;
	#10 counter$count = 74162;
	#10 counter$count = 74163;
	#10 counter$count = 74164;
	#10 counter$count = 74165;
	#10 counter$count = 74166;
	#10 counter$count = 74167;
	#10 counter$count = 74168;
	#10 counter$count = 74169;
	#10 counter$count = 74170;
	#10 counter$count = 74171;
	#10 counter$count = 74172;
	#10 counter$count = 74173;
	#10 counter$count = 74174;
	#10 counter$count = 74175;
	#10 counter$count = 74176;
	#10 counter$count = 74177;
	#10 counter$count = 74178;
	#10 counter$count = 74179;
	#10 counter$count = 74180;
	#10 counter$count = 74181;
	#10 counter$count = 74182;
	#10 counter$count = 74183;
	#10 counter$count = 74184;
	#10 counter$count = 74185;
	#10 counter$count = 74186;
	#10 counter$count = 74187;
	#10 counter$count = 74188;
	#10 counter$count = 74189;
	#10 counter$count = 74190;
	#10 counter$count = 74191;
	#10 counter$count = 74192;
	#10 counter$count = 74193;
	#10 counter$count = 74194;
	#10 counter$count = 74195;
	#10 counter$count = 74196;
	#10 counter$count = 74197;
	#10 counter$count = 74198;
	#10 counter$count = 74199;
	#10 counter$count = 74200;
	#10 counter$count = 74201;
	#10 counter$count = 74202;
	#10 counter$count = 74203;
	#10 counter$count = 74204;
	#10 counter$count = 74205;
	#10 counter$count = 74206;
	#10 counter$count = 74207;
	#10 counter$count = 74208;
	#10 counter$count = 74209;
	#10 counter$count = 74210;
	#10 counter$count = 74211;
	#10 counter$count = 74212;
	#10 counter$count = 74213;
	#10 counter$count = 74214;
	#10 counter$count = 74215;
	#10 counter$count = 74216;
	#10 counter$count = 74217;
	#10 counter$count = 74218;
	#10 counter$count = 74219;
	#10 counter$count = 74220;
	#10 counter$count = 74221;
	#10 counter$count = 74222;
	#10 counter$count = 74223;
	#10 counter$count = 74224;
	#10 counter$count = 74225;
	#10 counter$count = 74226;
	#10 counter$count = 74227;
	#10 counter$count = 74228;
	#10 counter$count = 74229;
	#10 counter$count = 74230;
	#10 counter$count = 74231;
	#10 counter$count = 74232;
	#10 counter$count = 74233;
	#10 counter$count = 74234;
	#10 counter$count = 74235;
	#10 counter$count = 74236;
	#10 counter$count = 74237;
	#10 counter$count = 74238;
	#10 counter$count = 74239;
	#10 counter$count = 74240;
	#10 counter$count = 74241;
	#10 counter$count = 74242;
	#10 counter$count = 74243;
	#10 counter$count = 74244;
	#10 counter$count = 74245;
	#10 counter$count = 74246;
	#10 counter$count = 74247;
	#10 counter$count = 74248;
	#10 counter$count = 74249;
	#10 counter$count = 74250;
	#10 counter$count = 74251;
	#10 counter$count = 74252;
	#10 counter$count = 74253;
	#10 counter$count = 74254;
	#10 counter$count = 74255;
	#10 counter$count = 74256;
	#10 counter$count = 74257;
	#10 counter$count = 74258;
	#10 counter$count = 74259;
	#10 counter$count = 74260;
	#10 counter$count = 74261;
	#10 counter$count = 74262;
	#10 counter$count = 74263;
	#10 counter$count = 74264;
	#10 counter$count = 74265;
	#10 counter$count = 74266;
	#10 counter$count = 74267;
	#10 counter$count = 74268;
	#10 counter$count = 74269;
	#10 counter$count = 74270;
	#10 counter$count = 74271;
	#10 counter$count = 74272;
	#10 counter$count = 74273;
	#10 counter$count = 74274;
	#10 counter$count = 74275;
	#10 counter$count = 74276;
	#10 counter$count = 74277;
	#10 counter$count = 74278;
	#10 counter$count = 74279;
	#10 counter$count = 74280;
	#10 counter$count = 74281;
	#10 counter$count = 74282;
	#10 counter$count = 74283;
	#10 counter$count = 74284;
	#10 counter$count = 74285;
	#10 counter$count = 74286;
	#10 counter$count = 74287;
	#10 counter$count = 74288;
	#10 counter$count = 74289;
	#10 counter$count = 74290;
	#10 counter$count = 74291;
	#10 counter$count = 74292;
	#10 counter$count = 74293;
	#10 counter$count = 74294;
	#10 counter$count = 74295;
	#10 counter$count = 74296;
	#10 counter$count = 74297;
	#10 counter$count = 74298;
	#10 counter$count = 74299;
	#10 counter$count = 74300;
	#10 counter$count = 74301;
	#10 counter$count = 74302;
	#10 counter$count = 74303;
	#10 counter$count = 74304;
	#10 counter$count = 74305;
	#10 counter$count = 74306;
	#10 counter$count = 74307;
	#10 counter$count = 74308;
	#10 counter$count = 74309;
	#10 counter$count = 74310;
	#10 counter$count = 74311;
	#10 counter$count = 74312;
	#10 counter$count = 74313;
	#10 counter$count = 74314;
	#10 counter$count = 74315;
	#10 counter$count = 74316;
	#10 counter$count = 74317;
	#10 counter$count = 74318;
	#10 counter$count = 74319;
	#10 counter$count = 74320;
	#10 counter$count = 74321;
	#10 counter$count = 74322;
	#10 counter$count = 74323;
	#10 counter$count = 74324;
	#10 counter$count = 74325;
	#10 counter$count = 74326;
	#10 counter$count = 74327;
	#10 counter$count = 74328;
	#10 counter$count = 74329;
	#10 counter$count = 74330;
	#10 counter$count = 74331;
	#10 counter$count = 74332;
	#10 counter$count = 74333;
	#10 counter$count = 74334;
	#10 counter$count = 74335;
	#10 counter$count = 74336;
	#10 counter$count = 74337;
	#10 counter$count = 74338;
	#10 counter$count = 74339;
	#10 counter$count = 74340;
	#10 counter$count = 74341;
	#10 counter$count = 74342;
	#10 counter$count = 74343;
	#10 counter$count = 74344;
	#10 counter$count = 74345;
	#10 counter$count = 74346;
	#10 counter$count = 74347;
	#10 counter$count = 74348;
	#10 counter$count = 74349;
	#10 counter$count = 74350;
	#10 counter$count = 74351;
	#10 counter$count = 74352;
	#10 counter$count = 74353;
	#10 counter$count = 74354;
	#10 counter$count = 74355;
	#10 counter$count = 74356;
	#10 counter$count = 74357;
	#10 counter$count = 74358;
	#10 counter$count = 74359;
	#10 counter$count = 74360;
	#10 counter$count = 74361;
	#10 counter$count = 74362;
	#10 counter$count = 74363;
	#10 counter$count = 74364;
	#10 counter$count = 74365;
	#10 counter$count = 74366;
	#10 counter$count = 74367;
	#10 counter$count = 74368;
	#10 counter$count = 74369;
	#10 counter$count = 74370;
	#10 counter$count = 74371;
	#10 counter$count = 74372;
	#10 counter$count = 74373;
	#10 counter$count = 74374;
	#10 counter$count = 74375;
	#10 counter$count = 74376;
	#10 counter$count = 74377;
	#10 counter$count = 74378;
	#10 counter$count = 74379;
	#10 counter$count = 74380;
	#10 counter$count = 74381;
	#10 counter$count = 74382;
	#10 counter$count = 74383;
	#10 counter$count = 74384;
	#10 counter$count = 74385;
	#10 counter$count = 74386;
	#10 counter$count = 74387;
	#10 counter$count = 74388;
	#10 counter$count = 74389;
	#10 counter$count = 74390;
	#10 counter$count = 74391;
	#10 counter$count = 74392;
	#10 counter$count = 74393;
	#10 counter$count = 74394;
	#10 counter$count = 74395;
	#10 counter$count = 74396;
	#10 counter$count = 74397;
	#10 counter$count = 74398;
	#10 counter$count = 74399;
	#10 counter$count = 74400;
	#10 counter$count = 74401;
	#10 counter$count = 74402;
	#10 counter$count = 74403;
	#10 counter$count = 74404;
	#10 counter$count = 74405;
	#10 counter$count = 74406;
	#10 counter$count = 74407;
	#10 counter$count = 74408;
	#10 counter$count = 74409;
	#10 counter$count = 74410;
	#10 counter$count = 74411;
	#10 counter$count = 74412;
	#10 counter$count = 74413;
	#10 counter$count = 74414;
	#10 counter$count = 74415;
	#10 counter$count = 74416;
	#10 counter$count = 74417;
	#10 counter$count = 74418;
	#10 counter$count = 74419;
	#10 counter$count = 74420;
	#10 counter$count = 74421;
	#10 counter$count = 74422;
	#10 counter$count = 74423;
	#10 counter$count = 74424;
	#10 counter$count = 74425;
	#10 counter$count = 74426;
	#10 counter$count = 74427;
	#10 counter$count = 74428;
	#10 counter$count = 74429;
	#10 counter$count = 74430;
	#10 counter$count = 74431;
	#10 counter$count = 74432;
	#10 counter$count = 74433;
	#10 counter$count = 74434;
	#10 counter$count = 74435;
	#10 counter$count = 74436;
	#10 counter$count = 74437;
	#10 counter$count = 74438;
	#10 counter$count = 74439;
	#10 counter$count = 74440;
	#10 counter$count = 74441;
	#10 counter$count = 74442;
	#10 counter$count = 74443;
	#10 counter$count = 74444;
	#10 counter$count = 74445;
	#10 counter$count = 74446;
	#10 counter$count = 74447;
	#10 counter$count = 74448;
	#10 counter$count = 74449;
	#10 counter$count = 74450;
	#10 counter$count = 74451;
	#10 counter$count = 74452;
	#10 counter$count = 74453;
	#10 counter$count = 74454;
	#10 counter$count = 74455;
	#10 counter$count = 74456;
	#10 counter$count = 74457;
	#10 counter$count = 74458;
	#10 counter$count = 74459;
	#10 counter$count = 74460;
	#10 counter$count = 74461;
	#10 counter$count = 74462;
	#10 counter$count = 74463;
	#10 counter$count = 74464;
	#10 counter$count = 74465;
	#10 counter$count = 74466;
	#10 counter$count = 74467;
	#10 counter$count = 74468;
	#10 counter$count = 74469;
	#10 counter$count = 74470;
	#10 counter$count = 74471;
	#10 counter$count = 74472;
	#10 counter$count = 74473;
	#10 counter$count = 74474;
	#10 counter$count = 74475;
	#10 counter$count = 74476;
	#10 counter$count = 74477;
	#10 counter$count = 74478;
	#10 counter$count = 74479;
	#10 counter$count = 74480;
	#10 counter$count = 74481;
	#10 counter$count = 74482;
	#10 counter$count = 74483;
	#10 counter$count = 74484;
	#10 counter$count = 74485;
	#10 counter$count = 74486;
	#10 counter$count = 74487;
	#10 counter$count = 74488;
	#10 counter$count = 74489;
	#10 counter$count = 74490;
	#10 counter$count = 74491;
	#10 counter$count = 74492;
	#10 counter$count = 74493;
	#10 counter$count = 74494;
	#10 counter$count = 74495;
	#10 counter$count = 74496;
	#10 counter$count = 74497;
	#10 counter$count = 74498;
	#10 counter$count = 74499;
	#10 counter$count = 74500;
	#10 counter$count = 74501;
	#10 counter$count = 74502;
	#10 counter$count = 74503;
	#10 counter$count = 74504;
	#10 counter$count = 74505;
	#10 counter$count = 74506;
	#10 counter$count = 74507;
	#10 counter$count = 74508;
	#10 counter$count = 74509;
	#10 counter$count = 74510;
	#10 counter$count = 74511;
	#10 counter$count = 74512;
	#10 counter$count = 74513;
	#10 counter$count = 74514;
	#10 counter$count = 74515;
	#10 counter$count = 74516;
	#10 counter$count = 74517;
	#10 counter$count = 74518;
	#10 counter$count = 74519;
	#10 counter$count = 74520;
	#10 counter$count = 74521;
	#10 counter$count = 74522;
	#10 counter$count = 74523;
	#10 counter$count = 74524;
	#10 counter$count = 74525;
	#10 counter$count = 74526;
	#10 counter$count = 74527;
	#10 counter$count = 74528;
	#10 counter$count = 74529;
	#10 counter$count = 74530;
	#10 counter$count = 74531;
	#10 counter$count = 74532;
	#10 counter$count = 74533;
	#10 counter$count = 74534;
	#10 counter$count = 74535;
	#10 counter$count = 74536;
	#10 counter$count = 74537;
	#10 counter$count = 74538;
	#10 counter$count = 74539;
	#10 counter$count = 74540;
	#10 counter$count = 74541;
	#10 counter$count = 74542;
	#10 counter$count = 74543;
	#10 counter$count = 74544;
	#10 counter$count = 74545;
	#10 counter$count = 74546;
	#10 counter$count = 74547;
	#10 counter$count = 74548;
	#10 counter$count = 74549;
	#10 counter$count = 74550;
	#10 counter$count = 74551;
	#10 counter$count = 74552;
	#10 counter$count = 74553;
	#10 counter$count = 74554;
	#10 counter$count = 74555;
	#10 counter$count = 74556;
	#10 counter$count = 74557;
	#10 counter$count = 74558;
	#10 counter$count = 74559;
	#10 counter$count = 74560;
	#10 counter$count = 74561;
	#10 counter$count = 74562;
	#10 counter$count = 74563;
	#10 counter$count = 74564;
	#10 counter$count = 74565;
	#10 counter$count = 74566;
	#10 counter$count = 74567;
	#10 counter$count = 74568;
	#10 counter$count = 74569;
	#10 counter$count = 74570;
	#10 counter$count = 74571;
	#10 counter$count = 74572;
	#10 counter$count = 74573;
	#10 counter$count = 74574;
	#10 counter$count = 74575;
	#10 counter$count = 74576;
	#10 counter$count = 74577;
	#10 counter$count = 74578;
	#10 counter$count = 74579;
	#10 counter$count = 74580;
	#10 counter$count = 74581;
	#10 counter$count = 74582;
	#10 counter$count = 74583;
	#10 counter$count = 74584;
	#10 counter$count = 74585;
	#10 counter$count = 74586;
	#10 counter$count = 74587;
	#10 counter$count = 74588;
	#10 counter$count = 74589;
	#10 counter$count = 74590;
	#10 counter$count = 74591;
	#10 counter$count = 74592;
	#10 counter$count = 74593;
	#10 counter$count = 74594;
	#10 counter$count = 74595;
	#10 counter$count = 74596;
	#10 counter$count = 74597;
	#10 counter$count = 74598;
	#10 counter$count = 74599;
	#10 counter$count = 74600;
	#10 counter$count = 74601;
	#10 counter$count = 74602;
	#10 counter$count = 74603;
	#10 counter$count = 74604;
	#10 counter$count = 74605;
	#10 counter$count = 74606;
	#10 counter$count = 74607;
	#10 counter$count = 74608;
	#10 counter$count = 74609;
	#10 counter$count = 74610;
	#10 counter$count = 74611;
	#10 counter$count = 74612;
	#10 counter$count = 74613;
	#10 counter$count = 74614;
	#10 counter$count = 74615;
	#10 counter$count = 74616;
	#10 counter$count = 74617;
	#10 counter$count = 74618;
	#10 counter$count = 74619;
	#10 counter$count = 74620;
	#10 counter$count = 74621;
	#10 counter$count = 74622;
	#10 counter$count = 74623;
	#10 counter$count = 74624;
	#10 counter$count = 74625;
	#10 counter$count = 74626;
	#10 counter$count = 74627;
	#10 counter$count = 74628;
	#10 counter$count = 74629;
	#10 counter$count = 74630;
	#10 counter$count = 74631;
	#10 counter$count = 74632;
	#10 counter$count = 74633;
	#10 counter$count = 74634;
	#10 counter$count = 74635;
	#10 counter$count = 74636;
	#10 counter$count = 74637;
	#10 counter$count = 74638;
	#10 counter$count = 74639;
	#10 counter$count = 74640;
	#10 counter$count = 74641;
	#10 counter$count = 74642;
	#10 counter$count = 74643;
	#10 counter$count = 74644;
	#10 counter$count = 74645;
	#10 counter$count = 74646;
	#10 counter$count = 74647;
	#10 counter$count = 74648;
	#10 counter$count = 74649;
	#10 counter$count = 74650;
	#10 counter$count = 74651;
	#10 counter$count = 74652;
	#10 counter$count = 74653;
	#10 counter$count = 74654;
	#10 counter$count = 74655;
	#10 counter$count = 74656;
	#10 counter$count = 74657;
	#10 counter$count = 74658;
	#10 counter$count = 74659;
	#10 counter$count = 74660;
	#10 counter$count = 74661;
	#10 counter$count = 74662;
	#10 counter$count = 74663;
	#10 counter$count = 74664;
	#10 counter$count = 74665;
	#10 counter$count = 74666;
	#10 counter$count = 74667;
	#10 counter$count = 74668;
	#10 counter$count = 74669;
	#10 counter$count = 74670;
	#10 counter$count = 74671;
	#10 counter$count = 74672;
	#10 counter$count = 74673;
	#10 counter$count = 74674;
	#10 counter$count = 74675;
	#10 counter$count = 74676;
	#10 counter$count = 74677;
	#10 counter$count = 74678;
	#10 counter$count = 74679;
	#10 counter$count = 74680;
	#10 counter$count = 74681;
	#10 counter$count = 74682;
	#10 counter$count = 74683;
	#10 counter$count = 74684;
	#10 counter$count = 74685;
	#10 counter$count = 74686;
	#10 counter$count = 74687;
	#10 counter$count = 74688;
	#10 counter$count = 74689;
	#10 counter$count = 74690;
	#10 counter$count = 74691;
	#10 counter$count = 74692;
	#10 counter$count = 74693;
	#10 counter$count = 74694;
	#10 counter$count = 74695;
	#10 counter$count = 74696;
	#10 counter$count = 74697;
	#10 counter$count = 74698;
	#10 counter$count = 74699;
	#10 counter$count = 74700;
	#10 counter$count = 74701;
	#10 counter$count = 74702;
	#10 counter$count = 74703;
	#10 counter$count = 74704;
	#10 counter$count = 74705;
	#10 counter$count = 74706;
	#10 counter$count = 74707;
	#10 counter$count = 74708;
	#10 counter$count = 74709;
	#10 counter$count = 74710;
	#10 counter$count = 74711;
	#10 counter$count = 74712;
	#10 counter$count = 74713;
	#10 counter$count = 74714;
	#10 counter$count = 74715;
	#10 counter$count = 74716;
	#10 counter$count = 74717;
	#10 counter$count = 74718;
	#10 counter$count = 74719;
	#10 counter$count = 74720;
	#10 counter$count = 74721;
	#10 counter$count = 74722;
	#10 counter$count = 74723;
	#10 counter$count = 74724;
	#10 counter$count = 74725;
	#10 counter$count = 74726;
	#10 counter$count = 74727;
	#10 counter$count = 74728;
	#10 counter$count = 74729;
	#10 counter$count = 74730;
	#10 counter$count = 74731;
	#10 counter$count = 74732;
	#10 counter$count = 74733;
	#10 counter$count = 74734;
	#10 counter$count = 74735;
	#10 counter$count = 74736;
	#10 counter$count = 74737;
	#10 counter$count = 74738;
	#10 counter$count = 74739;
	#10 counter$count = 74740;
	#10 counter$count = 74741;
	#10 counter$count = 74742;
	#10 counter$count = 74743;
	#10 counter$count = 74744;
	#10 counter$count = 74745;
	#10 counter$count = 74746;
	#10 counter$count = 74747;
	#10 counter$count = 74748;
	#10 counter$count = 74749;
	#10 counter$count = 74750;
	#10 counter$count = 74751;
	#10 counter$count = 74752;
	#10 counter$count = 74753;
	#10 counter$count = 74754;
	#10 counter$count = 74755;
	#10 counter$count = 74756;
	#10 counter$count = 74757;
	#10 counter$count = 74758;
	#10 counter$count = 74759;
	#10 counter$count = 74760;
	#10 counter$count = 74761;
	#10 counter$count = 74762;
	#10 counter$count = 74763;
	#10 counter$count = 74764;
	#10 counter$count = 74765;
	#10 counter$count = 74766;
	#10 counter$count = 74767;
	#10 counter$count = 74768;
	#10 counter$count = 74769;
	#10 counter$count = 74770;
	#10 counter$count = 74771;
	#10 counter$count = 74772;
	#10 counter$count = 74773;
	#10 counter$count = 74774;
	#10 counter$count = 74775;
	#10 counter$count = 74776;
	#10 counter$count = 74777;
	#10 counter$count = 74778;
	#10 counter$count = 74779;
	#10 counter$count = 74780;
	#10 counter$count = 74781;
	#10 counter$count = 74782;
	#10 counter$count = 74783;
	#10 counter$count = 74784;
	#10 counter$count = 74785;
	#10 counter$count = 74786;
	#10 counter$count = 74787;
	#10 counter$count = 74788;
	#10 counter$count = 74789;
	#10 counter$count = 74790;
	#10 counter$count = 74791;
	#10 counter$count = 74792;
	#10 counter$count = 74793;
	#10 counter$count = 74794;
	#10 counter$count = 74795;
	#10 counter$count = 74796;
	#10 counter$count = 74797;
	#10 counter$count = 74798;
	#10 counter$count = 74799;
	#10 counter$count = 74800;
	#10 counter$count = 74801;
	#10 counter$count = 74802;
	#10 counter$count = 74803;
	#10 counter$count = 74804;
	#10 counter$count = 74805;
	#10 counter$count = 74806;
	#10 counter$count = 74807;
	#10 counter$count = 74808;
	#10 counter$count = 74809;
	#10 counter$count = 74810;
	#10 counter$count = 74811;
	#10 counter$count = 74812;
	#10 counter$count = 74813;
	#10 counter$count = 74814;
	#10 counter$count = 74815;
	#10 counter$count = 74816;
	#10 counter$count = 74817;
	#10 counter$count = 74818;
	#10 counter$count = 74819;
	#10 counter$count = 74820;
	#10 counter$count = 74821;
	#10 counter$count = 74822;
	#10 counter$count = 74823;
	#10 counter$count = 74824;
	#10 counter$count = 74825;
	#10 counter$count = 74826;
	#10 counter$count = 74827;
	#10 counter$count = 74828;
	#10 counter$count = 74829;
	#10 counter$count = 74830;
	#10 counter$count = 74831;
	#10 counter$count = 74832;
	#10 counter$count = 74833;
	#10 counter$count = 74834;
	#10 counter$count = 74835;
	#10 counter$count = 74836;
	#10 counter$count = 74837;
	#10 counter$count = 74838;
	#10 counter$count = 74839;
	#10 counter$count = 74840;
	#10 counter$count = 74841;
	#10 counter$count = 74842;
	#10 counter$count = 74843;
	#10 counter$count = 74844;
	#10 counter$count = 74845;
	#10 counter$count = 74846;
	#10 counter$count = 74847;
	#10 counter$count = 74848;
	#10 counter$count = 74849;
	#10 counter$count = 74850;
	#10 counter$count = 74851;
	#10 counter$count = 74852;
	#10 counter$count = 74853;
	#10 counter$count = 74854;
	#10 counter$count = 74855;
	#10 counter$count = 74856;
	#10 counter$count = 74857;
	#10 counter$count = 74858;
	#10 counter$count = 74859;
	#10 counter$count = 74860;
	#10 counter$count = 74861;
	#10 counter$count = 74862;
	#10 counter$count = 74863;
	#10 counter$count = 74864;
	#10 counter$count = 74865;
	#10 counter$count = 74866;
	#10 counter$count = 74867;
	#10 counter$count = 74868;
	#10 counter$count = 74869;
	#10 counter$count = 74870;
	#10 counter$count = 74871;
	#10 counter$count = 74872;
	#10 counter$count = 74873;
	#10 counter$count = 74874;
	#10 counter$count = 74875;
	#10 counter$count = 74876;
	#10 counter$count = 74877;
	#10 counter$count = 74878;
	#10 counter$count = 74879;
	#10 counter$count = 74880;
	#10 counter$count = 74881;
	#10 counter$count = 74882;
	#10 counter$count = 74883;
	#10 counter$count = 74884;
	#10 counter$count = 74885;
	#10 counter$count = 74886;
	#10 counter$count = 74887;
	#10 counter$count = 74888;
	#10 counter$count = 74889;
	#10 counter$count = 74890;
	#10 counter$count = 74891;
	#10 counter$count = 74892;
	#10 counter$count = 74893;
	#10 counter$count = 74894;
	#10 counter$count = 74895;
	#10 counter$count = 74896;
	#10 counter$count = 74897;
	#10 counter$count = 74898;
	#10 counter$count = 74899;
	#10 counter$count = 74900;
	#10 counter$count = 74901;
	#10 counter$count = 74902;
	#10 counter$count = 74903;
	#10 counter$count = 74904;
	#10 counter$count = 74905;
	#10 counter$count = 74906;
	#10 counter$count = 74907;
	#10 counter$count = 74908;
	#10 counter$count = 74909;
	#10 counter$count = 74910;
	#10 counter$count = 74911;
	#10 counter$count = 74912;
	#10 counter$count = 74913;
	#10 counter$count = 74914;
	#10 counter$count = 74915;
	#10 counter$count = 74916;
	#10 counter$count = 74917;
	#10 counter$count = 74918;
	#10 counter$count = 74919;
	#10 counter$count = 74920;
	#10 counter$count = 74921;
	#10 counter$count = 74922;
	#10 counter$count = 74923;
	#10 counter$count = 74924;
	#10 counter$count = 74925;
	#10 counter$count = 74926;
	#10 counter$count = 74927;
	#10 counter$count = 74928;
	#10 counter$count = 74929;
	#10 counter$count = 74930;
	#10 counter$count = 74931;
	#10 counter$count = 74932;
	#10 counter$count = 74933;
	#10 counter$count = 74934;
	#10 counter$count = 74935;
	#10 counter$count = 74936;
	#10 counter$count = 74937;
	#10 counter$count = 74938;
	#10 counter$count = 74939;
	#10 counter$count = 74940;
	#10 counter$count = 74941;
	#10 counter$count = 74942;
	#10 counter$count = 74943;
	#10 counter$count = 74944;
	#10 counter$count = 74945;
	#10 counter$count = 74946;
	#10 counter$count = 74947;
	#10 counter$count = 74948;
	#10 counter$count = 74949;
	#10 counter$count = 74950;
	#10 counter$count = 74951;
	#10 counter$count = 74952;
	#10 counter$count = 74953;
	#10 counter$count = 74954;
	#10 counter$count = 74955;
	#10 counter$count = 74956;
	#10 counter$count = 74957;
	#10 counter$count = 74958;
	#10 counter$count = 74959;
	#10 counter$count = 74960;
	#10 counter$count = 74961;
	#10 counter$count = 74962;
	#10 counter$count = 74963;
	#10 counter$count = 74964;
	#10 counter$count = 74965;
	#10 counter$count = 74966;
	#10 counter$count = 74967;
	#10 counter$count = 74968;
	#10 counter$count = 74969;
	#10 counter$count = 74970;
	#10 counter$count = 74971;
	#10 counter$count = 74972;
	#10 counter$count = 74973;
	#10 counter$count = 74974;
	#10 counter$count = 74975;
	#10 counter$count = 74976;
	#10 counter$count = 74977;
	#10 counter$count = 74978;
	#10 counter$count = 74979;
	#10 counter$count = 74980;
	#10 counter$count = 74981;
	#10 counter$count = 74982;
	#10 counter$count = 74983;
	#10 counter$count = 74984;
	#10 counter$count = 74985;
	#10 counter$count = 74986;
	#10 counter$count = 74987;
	#10 counter$count = 74988;
	#10 counter$count = 74989;
	#10 counter$count = 74990;
	#10 counter$count = 74991;
	#10 counter$count = 74992;
	#10 counter$count = 74993;
	#10 counter$count = 74994;
	#10 counter$count = 74995;
	#10 counter$count = 74996;
	#10 counter$count = 74997;
	#10 counter$count = 74998;
	#10 counter$count = 74999;
	#10 counter$count = 75000;
	#10 counter$count = 75001;
	#10 counter$count = 75002;
	#10 counter$count = 75003;
	#10 counter$count = 75004;
	#10 counter$count = 75005;
	#10 counter$count = 75006;
	#10 counter$count = 75007;
	#10 counter$count = 75008;
	#10 counter$count = 75009;
	#10 counter$count = 75010;
	#10 counter$count = 75011;
	#10 counter$count = 75012;
	#10 counter$count = 75013;
	#10 counter$count = 75014;
	#10 counter$count = 75015;
	#10 counter$count = 75016;
	#10 counter$count = 75017;
	#10 counter$count = 75018;
	#10 counter$count = 75019;
	#10 counter$count = 75020;
	#10 counter$count = 75021;
	#10 counter$count = 75022;
	#10 counter$count = 75023;
	#10 counter$count = 75024;
	#10 counter$count = 75025;
	#10 counter$count = 75026;
	#10 counter$count = 75027;
	#10 counter$count = 75028;
	#10 counter$count = 75029;
	#10 counter$count = 75030;
	#10 counter$count = 75031;
	#10 counter$count = 75032;
	#10 counter$count = 75033;
	#10 counter$count = 75034;
	#10 counter$count = 75035;
	#10 counter$count = 75036;
	#10 counter$count = 75037;
	#10 counter$count = 75038;
	#10 counter$count = 75039;
	#10 counter$count = 75040;
	#10 counter$count = 75041;
	#10 counter$count = 75042;
	#10 counter$count = 75043;
	#10 counter$count = 75044;
	#10 counter$count = 75045;
	#10 counter$count = 75046;
	#10 counter$count = 75047;
	#10 counter$count = 75048;
	#10 counter$count = 75049;
	#10 counter$count = 75050;
	#10 counter$count = 75051;
	#10 counter$count = 75052;
	#10 counter$count = 75053;
	#10 counter$count = 75054;
	#10 counter$count = 75055;
	#10 counter$count = 75056;
	#10 counter$count = 75057;
	#10 counter$count = 75058;
	#10 counter$count = 75059;
	#10 counter$count = 75060;
	#10 counter$count = 75061;
	#10 counter$count = 75062;
	#10 counter$count = 75063;
	#10 counter$count = 75064;
	#10 counter$count = 75065;
	#10 counter$count = 75066;
	#10 counter$count = 75067;
	#10 counter$count = 75068;
	#10 counter$count = 75069;
	#10 counter$count = 75070;
	#10 counter$count = 75071;
	#10 counter$count = 75072;
	#10 counter$count = 75073;
	#10 counter$count = 75074;
	#10 counter$count = 75075;
	#10 counter$count = 75076;
	#10 counter$count = 75077;
	#10 counter$count = 75078;
	#10 counter$count = 75079;
	#10 counter$count = 75080;
	#10 counter$count = 75081;
	#10 counter$count = 75082;
	#10 counter$count = 75083;
	#10 counter$count = 75084;
	#10 counter$count = 75085;
	#10 counter$count = 75086;
	#10 counter$count = 75087;
	#10 counter$count = 75088;
	#10 counter$count = 75089;
	#10 counter$count = 75090;
	#10 counter$count = 75091;
	#10 counter$count = 75092;
	#10 counter$count = 75093;
	#10 counter$count = 75094;
	#10 counter$count = 75095;
	#10 counter$count = 75096;
	#10 counter$count = 75097;
	#10 counter$count = 75098;
	#10 counter$count = 75099;
	#10 counter$count = 75100;
	#10 counter$count = 75101;
	#10 counter$count = 75102;
	#10 counter$count = 75103;
	#10 counter$count = 75104;
	#10 counter$count = 75105;
	#10 counter$count = 75106;
	#10 counter$count = 75107;
	#10 counter$count = 75108;
	#10 counter$count = 75109;
	#10 counter$count = 75110;
	#10 counter$count = 75111;
	#10 counter$count = 75112;
	#10 counter$count = 75113;
	#10 counter$count = 75114;
	#10 counter$count = 75115;
	#10 counter$count = 75116;
	#10 counter$count = 75117;
	#10 counter$count = 75118;
	#10 counter$count = 75119;
	#10 counter$count = 75120;
	#10 counter$count = 75121;
	#10 counter$count = 75122;
	#10 counter$count = 75123;
	#10 counter$count = 75124;
	#10 counter$count = 75125;
	#10 counter$count = 75126;
	#10 counter$count = 75127;
	#10 counter$count = 75128;
	#10 counter$count = 75129;
	#10 counter$count = 75130;
	#10 counter$count = 75131;
	#10 counter$count = 75132;
	#10 counter$count = 75133;
	#10 counter$count = 75134;
	#10 counter$count = 75135;
	#10 counter$count = 75136;
	#10 counter$count = 75137;
	#10 counter$count = 75138;
	#10 counter$count = 75139;
	#10 counter$count = 75140;
	#10 counter$count = 75141;
	#10 counter$count = 75142;
	#10 counter$count = 75143;
	#10 counter$count = 75144;
	#10 counter$count = 75145;
	#10 counter$count = 75146;
	#10 counter$count = 75147;
	#10 counter$count = 75148;
	#10 counter$count = 75149;
	#10 counter$count = 75150;
	#10 counter$count = 75151;
	#10 counter$count = 75152;
	#10 counter$count = 75153;
	#10 counter$count = 75154;
	#10 counter$count = 75155;
	#10 counter$count = 75156;
	#10 counter$count = 75157;
	#10 counter$count = 75158;
	#10 counter$count = 75159;
	#10 counter$count = 75160;
	#10 counter$count = 75161;
	#10 counter$count = 75162;
	#10 counter$count = 75163;
	#10 counter$count = 75164;
	#10 counter$count = 75165;
	#10 counter$count = 75166;
	#10 counter$count = 75167;
	#10 counter$count = 75168;
	#10 counter$count = 75169;
	#10 counter$count = 75170;
	#10 counter$count = 75171;
	#10 counter$count = 75172;
	#10 counter$count = 75173;
	#10 counter$count = 75174;
	#10 counter$count = 75175;
	#10 counter$count = 75176;
	#10 counter$count = 75177;
	#10 counter$count = 75178;
	#10 counter$count = 75179;
	#10 counter$count = 75180;
	#10 counter$count = 75181;
	#10 counter$count = 75182;
	#10 counter$count = 75183;
	#10 counter$count = 75184;
	#10 counter$count = 75185;
	#10 counter$count = 75186;
	#10 counter$count = 75187;
	#10 counter$count = 75188;
	#10 counter$count = 75189;
	#10 counter$count = 75190;
	#10 counter$count = 75191;
	#10 counter$count = 75192;
	#10 counter$count = 75193;
	#10 counter$count = 75194;
	#10 counter$count = 75195;
	#10 counter$count = 75196;
	#10 counter$count = 75197;
	#10 counter$count = 75198;
	#10 counter$count = 75199;
	#10 counter$count = 75200;
	#10 counter$count = 75201;
	#10 counter$count = 75202;
	#10 counter$count = 75203;
	#10 counter$count = 75204;
	#10 counter$count = 75205;
	#10 counter$count = 75206;
	#10 counter$count = 75207;
	#10 counter$count = 75208;
	#10 counter$count = 75209;
	#10 counter$count = 75210;
	#10 counter$count = 75211;
	#10 counter$count = 75212;
	#10 counter$count = 75213;
	#10 counter$count = 75214;
	#10 counter$count = 75215;
	#10 counter$count = 75216;
	#10 counter$count = 75217;
	#10 counter$count = 75218;
	#10 counter$count = 75219;
	#10 counter$count = 75220;
	#10 counter$count = 75221;
	#10 counter$count = 75222;
	#10 counter$count = 75223;
	#10 counter$count = 75224;
	#10 counter$count = 75225;
	#10 counter$count = 75226;
	#10 counter$count = 75227;
	#10 counter$count = 75228;
	#10 counter$count = 75229;
	#10 counter$count = 75230;
	#10 counter$count = 75231;
	#10 counter$count = 75232;
	#10 counter$count = 75233;
	#10 counter$count = 75234;
	#10 counter$count = 75235;
	#10 counter$count = 75236;
	#10 counter$count = 75237;
	#10 counter$count = 75238;
	#10 counter$count = 75239;
	#10 counter$count = 75240;
	#10 counter$count = 75241;
	#10 counter$count = 75242;
	#10 counter$count = 75243;
	#10 counter$count = 75244;
	#10 counter$count = 75245;
	#10 counter$count = 75246;
	#10 counter$count = 75247;
	#10 counter$count = 75248;
	#10 counter$count = 75249;
	#10 counter$count = 75250;
	#10 counter$count = 75251;
	#10 counter$count = 75252;
	#10 counter$count = 75253;
	#10 counter$count = 75254;
	#10 counter$count = 75255;
	#10 counter$count = 75256;
	#10 counter$count = 75257;
	#10 counter$count = 75258;
	#10 counter$count = 75259;
	#10 counter$count = 75260;
	#10 counter$count = 75261;
	#10 counter$count = 75262;
	#10 counter$count = 75263;
	#10 counter$count = 75264;
	#10 counter$count = 75265;
	#10 counter$count = 75266;
	#10 counter$count = 75267;
	#10 counter$count = 75268;
	#10 counter$count = 75269;
	#10 counter$count = 75270;
	#10 counter$count = 75271;
	#10 counter$count = 75272;
	#10 counter$count = 75273;
	#10 counter$count = 75274;
	#10 counter$count = 75275;
	#10 counter$count = 75276;
	#10 counter$count = 75277;
	#10 counter$count = 75278;
	#10 counter$count = 75279;
	#10 counter$count = 75280;
	#10 counter$count = 75281;
	#10 counter$count = 75282;
	#10 counter$count = 75283;
	#10 counter$count = 75284;
	#10 counter$count = 75285;
	#10 counter$count = 75286;
	#10 counter$count = 75287;
	#10 counter$count = 75288;
	#10 counter$count = 75289;
	#10 counter$count = 75290;
	#10 counter$count = 75291;
	#10 counter$count = 75292;
	#10 counter$count = 75293;
	#10 counter$count = 75294;
	#10 counter$count = 75295;
	#10 counter$count = 75296;
	#10 counter$count = 75297;
	#10 counter$count = 75298;
	#10 counter$count = 75299;
	#10 counter$count = 75300;
	#10 counter$count = 75301;
	#10 counter$count = 75302;
	#10 counter$count = 75303;
	#10 counter$count = 75304;
	#10 counter$count = 75305;
	#10 counter$count = 75306;
	#10 counter$count = 75307;
	#10 counter$count = 75308;
	#10 counter$count = 75309;
	#10 counter$count = 75310;
	#10 counter$count = 75311;
	#10 counter$count = 75312;
	#10 counter$count = 75313;
	#10 counter$count = 75314;
	#10 counter$count = 75315;
	#10 counter$count = 75316;
	#10 counter$count = 75317;
	#10 counter$count = 75318;
	#10 counter$count = 75319;
	#10 counter$count = 75320;
	#10 counter$count = 75321;
	#10 counter$count = 75322;
	#10 counter$count = 75323;
	#10 counter$count = 75324;
	#10 counter$count = 75325;
	#10 counter$count = 75326;
	#10 counter$count = 75327;
	#10 counter$count = 75328;
	#10 counter$count = 75329;
	#10 counter$count = 75330;
	#10 counter$count = 75331;
	#10 counter$count = 75332;
	#10 counter$count = 75333;
	#10 counter$count = 75334;
	#10 counter$count = 75335;
	#10 counter$count = 75336;
	#10 counter$count = 75337;
	#10 counter$count = 75338;
	#10 counter$count = 75339;
	#10 counter$count = 75340;
	#10 counter$count = 75341;
	#10 counter$count = 75342;
	#10 counter$count = 75343;
	#10 counter$count = 75344;
	#10 counter$count = 75345;
	#10 counter$count = 75346;
	#10 counter$count = 75347;
	#10 counter$count = 75348;
	#10 counter$count = 75349;
	#10 counter$count = 75350;
	#10 counter$count = 75351;
	#10 counter$count = 75352;
	#10 counter$count = 75353;
	#10 counter$count = 75354;
	#10 counter$count = 75355;
	#10 counter$count = 75356;
	#10 counter$count = 75357;
	#10 counter$count = 75358;
	#10 counter$count = 75359;
	#10 counter$count = 75360;
	#10 counter$count = 75361;
	#10 counter$count = 75362;
	#10 counter$count = 75363;
	#10 counter$count = 75364;
	#10 counter$count = 75365;
	#10 counter$count = 75366;
	#10 counter$count = 75367;
	#10 counter$count = 75368;
	#10 counter$count = 75369;
	#10 counter$count = 75370;
	#10 counter$count = 75371;
	#10 counter$count = 75372;
	#10 counter$count = 75373;
	#10 counter$count = 75374;
	#10 counter$count = 75375;
	#10 counter$count = 75376;
	#10 counter$count = 75377;
	#10 counter$count = 75378;
	#10 counter$count = 75379;
	#10 counter$count = 75380;
	#10 counter$count = 75381;
	#10 counter$count = 75382;
	#10 counter$count = 75383;
	#10 counter$count = 75384;
	#10 counter$count = 75385;
	#10 counter$count = 75386;
	#10 counter$count = 75387;
	#10 counter$count = 75388;
	#10 counter$count = 75389;
	#10 counter$count = 75390;
	#10 counter$count = 75391;
	#10 counter$count = 75392;
	#10 counter$count = 75393;
	#10 counter$count = 75394;
	#10 counter$count = 75395;
	#10 counter$count = 75396;
	#10 counter$count = 75397;
	#10 counter$count = 75398;
	#10 counter$count = 75399;
	#10 counter$count = 75400;
	#10 counter$count = 75401;
	#10 counter$count = 75402;
	#10 counter$count = 75403;
	#10 counter$count = 75404;
	#10 counter$count = 75405;
	#10 counter$count = 75406;
	#10 counter$count = 75407;
	#10 counter$count = 75408;
	#10 counter$count = 75409;
	#10 counter$count = 75410;
	#10 counter$count = 75411;
	#10 counter$count = 75412;
	#10 counter$count = 75413;
	#10 counter$count = 75414;
	#10 counter$count = 75415;
	#10 counter$count = 75416;
	#10 counter$count = 75417;
	#10 counter$count = 75418;
	#10 counter$count = 75419;
	#10 counter$count = 75420;
	#10 counter$count = 75421;
	#10 counter$count = 75422;
	#10 counter$count = 75423;
	#10 counter$count = 75424;
	#10 counter$count = 75425;
	#10 counter$count = 75426;
	#10 counter$count = 75427;
	#10 counter$count = 75428;
	#10 counter$count = 75429;
	#10 counter$count = 75430;
	#10 counter$count = 75431;
	#10 counter$count = 75432;
	#10 counter$count = 75433;
	#10 counter$count = 75434;
	#10 counter$count = 75435;
	#10 counter$count = 75436;
	#10 counter$count = 75437;
	#10 counter$count = 75438;
	#10 counter$count = 75439;
	#10 counter$count = 75440;
	#10 counter$count = 75441;
	#10 counter$count = 75442;
	#10 counter$count = 75443;
	#10 counter$count = 75444;
	#10 counter$count = 75445;
	#10 counter$count = 75446;
	#10 counter$count = 75447;
	#10 counter$count = 75448;
	#10 counter$count = 75449;
	#10 counter$count = 75450;
	#10 counter$count = 75451;
	#10 counter$count = 75452;
	#10 counter$count = 75453;
	#10 counter$count = 75454;
	#10 counter$count = 75455;
	#10 counter$count = 75456;
	#10 counter$count = 75457;
	#10 counter$count = 75458;
	#10 counter$count = 75459;
	#10 counter$count = 75460;
	#10 counter$count = 75461;
	#10 counter$count = 75462;
	#10 counter$count = 75463;
	#10 counter$count = 75464;
	#10 counter$count = 75465;
	#10 counter$count = 75466;
	#10 counter$count = 75467;
	#10 counter$count = 75468;
	#10 counter$count = 75469;
	#10 counter$count = 75470;
	#10 counter$count = 75471;
	#10 counter$count = 75472;
	#10 counter$count = 75473;
	#10 counter$count = 75474;
	#10 counter$count = 75475;
	#10 counter$count = 75476;
	#10 counter$count = 75477;
	#10 counter$count = 75478;
	#10 counter$count = 75479;
	#10 counter$count = 75480;
	#10 counter$count = 75481;
	#10 counter$count = 75482;
	#10 counter$count = 75483;
	#10 counter$count = 75484;
	#10 counter$count = 75485;
	#10 counter$count = 75486;
	#10 counter$count = 75487;
	#10 counter$count = 75488;
	#10 counter$count = 75489;
	#10 counter$count = 75490;
	#10 counter$count = 75491;
	#10 counter$count = 75492;
	#10 counter$count = 75493;
	#10 counter$count = 75494;
	#10 counter$count = 75495;
	#10 counter$count = 75496;
	#10 counter$count = 75497;
	#10 counter$count = 75498;
	#10 counter$count = 75499;
	#10 counter$count = 75500;
	#10 counter$count = 75501;
	#10 counter$count = 75502;
	#10 counter$count = 75503;
	#10 counter$count = 75504;
	#10 counter$count = 75505;
	#10 counter$count = 75506;
	#10 counter$count = 75507;
	#10 counter$count = 75508;
	#10 counter$count = 75509;
	#10 counter$count = 75510;
	#10 counter$count = 75511;
	#10 counter$count = 75512;
	#10 counter$count = 75513;
	#10 counter$count = 75514;
	#10 counter$count = 75515;
	#10 counter$count = 75516;
	#10 counter$count = 75517;
	#10 counter$count = 75518;
	#10 counter$count = 75519;
	#10 counter$count = 75520;
	#10 counter$count = 75521;
	#10 counter$count = 75522;
	#10 counter$count = 75523;
	#10 counter$count = 75524;
	#10 counter$count = 75525;
	#10 counter$count = 75526;
	#10 counter$count = 75527;
	#10 counter$count = 75528;
	#10 counter$count = 75529;
	#10 counter$count = 75530;
	#10 counter$count = 75531;
	#10 counter$count = 75532;
	#10 counter$count = 75533;
	#10 counter$count = 75534;
	#10 counter$count = 75535;
	#10 counter$count = 75536;
	#10 counter$count = 75537;
	#10 counter$count = 75538;
	#10 counter$count = 75539;
	#10 counter$count = 75540;
	#10 counter$count = 75541;
	#10 counter$count = 75542;
	#10 counter$count = 75543;
	#10 counter$count = 75544;
	#10 counter$count = 75545;
	#10 counter$count = 75546;
	#10 counter$count = 75547;
	#10 counter$count = 75548;
	#10 counter$count = 75549;
	#10 counter$count = 75550;
	#10 counter$count = 75551;
	#10 counter$count = 75552;
	#10 counter$count = 75553;
	#10 counter$count = 75554;
	#10 counter$count = 75555;
	#10 counter$count = 75556;
	#10 counter$count = 75557;
	#10 counter$count = 75558;
	#10 counter$count = 75559;
	#10 counter$count = 75560;
	#10 counter$count = 75561;
	#10 counter$count = 75562;
	#10 counter$count = 75563;
	#10 counter$count = 75564;
	#10 counter$count = 75565;
	#10 counter$count = 75566;
	#10 counter$count = 75567;
	#10 counter$count = 75568;
	#10 counter$count = 75569;
	#10 counter$count = 75570;
	#10 counter$count = 75571;
	#10 counter$count = 75572;
	#10 counter$count = 75573;
	#10 counter$count = 75574;
	#10 counter$count = 75575;
	#10 counter$count = 75576;
	#10 counter$count = 75577;
	#10 counter$count = 75578;
	#10 counter$count = 75579;
	#10 counter$count = 75580;
	#10 counter$count = 75581;
	#10 counter$count = 75582;
	#10 counter$count = 75583;
	#10 counter$count = 75584;
	#10 counter$count = 75585;
	#10 counter$count = 75586;
	#10 counter$count = 75587;
	#10 counter$count = 75588;
	#10 counter$count = 75589;
	#10 counter$count = 75590;
	#10 counter$count = 75591;
	#10 counter$count = 75592;
	#10 counter$count = 75593;
	#10 counter$count = 75594;
	#10 counter$count = 75595;
	#10 counter$count = 75596;
	#10 counter$count = 75597;
	#10 counter$count = 75598;
	#10 counter$count = 75599;
	#10 counter$count = 75600;
	#10 counter$count = 75601;
	#10 counter$count = 75602;
	#10 counter$count = 75603;
	#10 counter$count = 75604;
	#10 counter$count = 75605;
	#10 counter$count = 75606;
	#10 counter$count = 75607;
	#10 counter$count = 75608;
	#10 counter$count = 75609;
	#10 counter$count = 75610;
	#10 counter$count = 75611;
	#10 counter$count = 75612;
	#10 counter$count = 75613;
	#10 counter$count = 75614;
	#10 counter$count = 75615;
	#10 counter$count = 75616;
	#10 counter$count = 75617;
	#10 counter$count = 75618;
	#10 counter$count = 75619;
	#10 counter$count = 75620;
	#10 counter$count = 75621;
	#10 counter$count = 75622;
	#10 counter$count = 75623;
	#10 counter$count = 75624;
	#10 counter$count = 75625;
	#10 counter$count = 75626;
	#10 counter$count = 75627;
	#10 counter$count = 75628;
	#10 counter$count = 75629;
	#10 counter$count = 75630;
	#10 counter$count = 75631;
	#10 counter$count = 75632;
	#10 counter$count = 75633;
	#10 counter$count = 75634;
	#10 counter$count = 75635;
	#10 counter$count = 75636;
	#10 counter$count = 75637;
	#10 counter$count = 75638;
	#10 counter$count = 75639;
	#10 counter$count = 75640;
	#10 counter$count = 75641;
	#10 counter$count = 75642;
	#10 counter$count = 75643;
	#10 counter$count = 75644;
	#10 counter$count = 75645;
	#10 counter$count = 75646;
	#10 counter$count = 75647;
	#10 counter$count = 75648;
	#10 counter$count = 75649;
	#10 counter$count = 75650;
	#10 counter$count = 75651;
	#10 counter$count = 75652;
	#10 counter$count = 75653;
	#10 counter$count = 75654;
	#10 counter$count = 75655;
	#10 counter$count = 75656;
	#10 counter$count = 75657;
	#10 counter$count = 75658;
	#10 counter$count = 75659;
	#10 counter$count = 75660;
	#10 counter$count = 75661;
	#10 counter$count = 75662;
	#10 counter$count = 75663;
	#10 counter$count = 75664;
	#10 counter$count = 75665;
	#10 counter$count = 75666;
	#10 counter$count = 75667;
	#10 counter$count = 75668;
	#10 counter$count = 75669;
	#10 counter$count = 75670;
	#10 counter$count = 75671;
	#10 counter$count = 75672;
	#10 counter$count = 75673;
	#10 counter$count = 75674;
	#10 counter$count = 75675;
	#10 counter$count = 75676;
	#10 counter$count = 75677;
	#10 counter$count = 75678;
	#10 counter$count = 75679;
	#10 counter$count = 75680;
	#10 counter$count = 75681;
	#10 counter$count = 75682;
	#10 counter$count = 75683;
	#10 counter$count = 75684;
	#10 counter$count = 75685;
	#10 counter$count = 75686;
	#10 counter$count = 75687;
	#10 counter$count = 75688;
	#10 counter$count = 75689;
	#10 counter$count = 75690;
	#10 counter$count = 75691;
	#10 counter$count = 75692;
	#10 counter$count = 75693;
	#10 counter$count = 75694;
	#10 counter$count = 75695;
	#10 counter$count = 75696;
	#10 counter$count = 75697;
	#10 counter$count = 75698;
	#10 counter$count = 75699;
	#10 counter$count = 75700;
	#10 counter$count = 75701;
	#10 counter$count = 75702;
	#10 counter$count = 75703;
	#10 counter$count = 75704;
	#10 counter$count = 75705;
	#10 counter$count = 75706;
	#10 counter$count = 75707;
	#10 counter$count = 75708;
	#10 counter$count = 75709;
	#10 counter$count = 75710;
	#10 counter$count = 75711;
	#10 counter$count = 75712;
	#10 counter$count = 75713;
	#10 counter$count = 75714;
	#10 counter$count = 75715;
	#10 counter$count = 75716;
	#10 counter$count = 75717;
	#10 counter$count = 75718;
	#10 counter$count = 75719;
	#10 counter$count = 75720;
	#10 counter$count = 75721;
	#10 counter$count = 75722;
	#10 counter$count = 75723;
	#10 counter$count = 75724;
	#10 counter$count = 75725;
	#10 counter$count = 75726;
	#10 counter$count = 75727;
	#10 counter$count = 75728;
	#10 counter$count = 75729;
	#10 counter$count = 75730;
	#10 counter$count = 75731;
	#10 counter$count = 75732;
	#10 counter$count = 75733;
	#10 counter$count = 75734;
	#10 counter$count = 75735;
	#10 counter$count = 75736;
	#10 counter$count = 75737;
	#10 counter$count = 75738;
	#10 counter$count = 75739;
	#10 counter$count = 75740;
	#10 counter$count = 75741;
	#10 counter$count = 75742;
	#10 counter$count = 75743;
	#10 counter$count = 75744;
	#10 counter$count = 75745;
	#10 counter$count = 75746;
	#10 counter$count = 75747;
	#10 counter$count = 75748;
	#10 counter$count = 75749;
	#10 counter$count = 75750;
	#10 counter$count = 75751;
	#10 counter$count = 75752;
	#10 counter$count = 75753;
	#10 counter$count = 75754;
	#10 counter$count = 75755;
	#10 counter$count = 75756;
	#10 counter$count = 75757;
	#10 counter$count = 75758;
	#10 counter$count = 75759;
	#10 counter$count = 75760;
	#10 counter$count = 75761;
	#10 counter$count = 75762;
	#10 counter$count = 75763;
	#10 counter$count = 75764;
	#10 counter$count = 75765;
	#10 counter$count = 75766;
	#10 counter$count = 75767;
	#10 counter$count = 75768;
	#10 counter$count = 75769;
	#10 counter$count = 75770;
	#10 counter$count = 75771;
	#10 counter$count = 75772;
	#10 counter$count = 75773;
	#10 counter$count = 75774;
	#10 counter$count = 75775;
	#10 counter$count = 75776;
	#10 counter$count = 75777;
	#10 counter$count = 75778;
	#10 counter$count = 75779;
	#10 counter$count = 75780;
	#10 counter$count = 75781;
	#10 counter$count = 75782;
	#10 counter$count = 75783;
	#10 counter$count = 75784;
	#10 counter$count = 75785;
	#10 counter$count = 75786;
	#10 counter$count = 75787;
	#10 counter$count = 75788;
	#10 counter$count = 75789;
	#10 counter$count = 75790;
	#10 counter$count = 75791;
	#10 counter$count = 75792;
	#10 counter$count = 75793;
	#10 counter$count = 75794;
	#10 counter$count = 75795;
	#10 counter$count = 75796;
	#10 counter$count = 75797;
	#10 counter$count = 75798;
	#10 counter$count = 75799;
	#10 counter$count = 75800;
	#10 counter$count = 75801;
	#10 counter$count = 75802;
	#10 counter$count = 75803;
	#10 counter$count = 75804;
	#10 counter$count = 75805;
	#10 counter$count = 75806;
	#10 counter$count = 75807;
	#10 counter$count = 75808;
	#10 counter$count = 75809;
	#10 counter$count = 75810;
	#10 counter$count = 75811;
	#10 counter$count = 75812;
	#10 counter$count = 75813;
	#10 counter$count = 75814;
	#10 counter$count = 75815;
	#10 counter$count = 75816;
	#10 counter$count = 75817;
	#10 counter$count = 75818;
	#10 counter$count = 75819;
	#10 counter$count = 75820;
	#10 counter$count = 75821;
	#10 counter$count = 75822;
	#10 counter$count = 75823;
	#10 counter$count = 75824;
	#10 counter$count = 75825;
	#10 counter$count = 75826;
	#10 counter$count = 75827;
	#10 counter$count = 75828;
	#10 counter$count = 75829;
	#10 counter$count = 75830;
	#10 counter$count = 75831;
	#10 counter$count = 75832;
	#10 counter$count = 75833;
	#10 counter$count = 75834;
	#10 counter$count = 75835;
	#10 counter$count = 75836;
	#10 counter$count = 75837;
	#10 counter$count = 75838;
	#10 counter$count = 75839;
	#10 counter$count = 75840;
	#10 counter$count = 75841;
	#10 counter$count = 75842;
	#10 counter$count = 75843;
	#10 counter$count = 75844;
	#10 counter$count = 75845;
	#10 counter$count = 75846;
	#10 counter$count = 75847;
	#10 counter$count = 75848;
	#10 counter$count = 75849;
	#10 counter$count = 75850;
	#10 counter$count = 75851;
	#10 counter$count = 75852;
	#10 counter$count = 75853;
	#10 counter$count = 75854;
	#10 counter$count = 75855;
	#10 counter$count = 75856;
	#10 counter$count = 75857;
	#10 counter$count = 75858;
	#10 counter$count = 75859;
	#10 counter$count = 75860;
	#10 counter$count = 75861;
	#10 counter$count = 75862;
	#10 counter$count = 75863;
	#10 counter$count = 75864;
	#10 counter$count = 75865;
	#10 counter$count = 75866;
	#10 counter$count = 75867;
	#10 counter$count = 75868;
	#10 counter$count = 75869;
	#10 counter$count = 75870;
	#10 counter$count = 75871;
	#10 counter$count = 75872;
	#10 counter$count = 75873;
	#10 counter$count = 75874;
	#10 counter$count = 75875;
	#10 counter$count = 75876;
	#10 counter$count = 75877;
	#10 counter$count = 75878;
	#10 counter$count = 75879;
	#10 counter$count = 75880;
	#10 counter$count = 75881;
	#10 counter$count = 75882;
	#10 counter$count = 75883;
	#10 counter$count = 75884;
	#10 counter$count = 75885;
	#10 counter$count = 75886;
	#10 counter$count = 75887;
	#10 counter$count = 75888;
	#10 counter$count = 75889;
	#10 counter$count = 75890;
	#10 counter$count = 75891;
	#10 counter$count = 75892;
	#10 counter$count = 75893;
	#10 counter$count = 75894;
	#10 counter$count = 75895;
	#10 counter$count = 75896;
	#10 counter$count = 75897;
	#10 counter$count = 75898;
	#10 counter$count = 75899;
	#10 counter$count = 75900;
	#10 counter$count = 75901;
	#10 counter$count = 75902;
	#10 counter$count = 75903;
	#10 counter$count = 75904;
	#10 counter$count = 75905;
	#10 counter$count = 75906;
	#10 counter$count = 75907;
	#10 counter$count = 75908;
	#10 counter$count = 75909;
	#10 counter$count = 75910;
	#10 counter$count = 75911;
	#10 counter$count = 75912;
	#10 counter$count = 75913;
	#10 counter$count = 75914;
	#10 counter$count = 75915;
	#10 counter$count = 75916;
	#10 counter$count = 75917;
	#10 counter$count = 75918;
	#10 counter$count = 75919;
	#10 counter$count = 75920;
	#10 counter$count = 75921;
	#10 counter$count = 75922;
	#10 counter$count = 75923;
	#10 counter$count = 75924;
	#10 counter$count = 75925;
	#10 counter$count = 75926;
	#10 counter$count = 75927;
	#10 counter$count = 75928;
	#10 counter$count = 75929;
	#10 counter$count = 75930;
	#10 counter$count = 75931;
	#10 counter$count = 75932;
	#10 counter$count = 75933;
	#10 counter$count = 75934;
	#10 counter$count = 75935;
	#10 counter$count = 75936;
	#10 counter$count = 75937;
	#10 counter$count = 75938;
	#10 counter$count = 75939;
	#10 counter$count = 75940;
	#10 counter$count = 75941;
	#10 counter$count = 75942;
	#10 counter$count = 75943;
	#10 counter$count = 75944;
	#10 counter$count = 75945;
	#10 counter$count = 75946;
	#10 counter$count = 75947;
	#10 counter$count = 75948;
	#10 counter$count = 75949;
	#10 counter$count = 75950;
	#10 counter$count = 75951;
	#10 counter$count = 75952;
	#10 counter$count = 75953;
	#10 counter$count = 75954;
	#10 counter$count = 75955;
	#10 counter$count = 75956;
	#10 counter$count = 75957;
	#10 counter$count = 75958;
	#10 counter$count = 75959;
	#10 counter$count = 75960;
	#10 counter$count = 75961;
	#10 counter$count = 75962;
	#10 counter$count = 75963;
	#10 counter$count = 75964;
	#10 counter$count = 75965;
	#10 counter$count = 75966;
	#10 counter$count = 75967;
	#10 counter$count = 75968;
	#10 counter$count = 75969;
	#10 counter$count = 75970;
	#10 counter$count = 75971;
	#10 counter$count = 75972;
	#10 counter$count = 75973;
	#10 counter$count = 75974;
	#10 counter$count = 75975;
	#10 counter$count = 75976;
	#10 counter$count = 75977;
	#10 counter$count = 75978;
	#10 counter$count = 75979;
	#10 counter$count = 75980;
	#10 counter$count = 75981;
	#10 counter$count = 75982;
	#10 counter$count = 75983;
	#10 counter$count = 75984;
	#10 counter$count = 75985;
	#10 counter$count = 75986;
	#10 counter$count = 75987;
	#10 counter$count = 75988;
	#10 counter$count = 75989;
	#10 counter$count = 75990;
	#10 counter$count = 75991;
	#10 counter$count = 75992;
	#10 counter$count = 75993;
	#10 counter$count = 75994;
	#10 counter$count = 75995;
	#10 counter$count = 75996;
	#10 counter$count = 75997;
	#10 counter$count = 75998;
	#10 counter$count = 75999;
	#10 counter$count = 76000;
	#10 counter$count = 76001;
	#10 counter$count = 76002;
	#10 counter$count = 76003;
	#10 counter$count = 76004;
	#10 counter$count = 76005;
	#10 counter$count = 76006;
	#10 counter$count = 76007;
	#10 counter$count = 76008;
	#10 counter$count = 76009;
	#10 counter$count = 76010;
	#10 counter$count = 76011;
	#10 counter$count = 76012;
	#10 counter$count = 76013;
	#10 counter$count = 76014;
	#10 counter$count = 76015;
	#10 counter$count = 76016;
	#10 counter$count = 76017;
	#10 counter$count = 76018;
	#10 counter$count = 76019;
	#10 counter$count = 76020;
	#10 counter$count = 76021;
	#10 counter$count = 76022;
	#10 counter$count = 76023;
	#10 counter$count = 76024;
	#10 counter$count = 76025;
	#10 counter$count = 76026;
	#10 counter$count = 76027;
	#10 counter$count = 76028;
	#10 counter$count = 76029;
	#10 counter$count = 76030;
	#10 counter$count = 76031;
	#10 counter$count = 76032;
	#10 counter$count = 76033;
	#10 counter$count = 76034;
	#10 counter$count = 76035;
	#10 counter$count = 76036;
	#10 counter$count = 76037;
	#10 counter$count = 76038;
	#10 counter$count = 76039;
	#10 counter$count = 76040;
	#10 counter$count = 76041;
	#10 counter$count = 76042;
	#10 counter$count = 76043;
	#10 counter$count = 76044;
	#10 counter$count = 76045;
	#10 counter$count = 76046;
	#10 counter$count = 76047;
	#10 counter$count = 76048;
	#10 counter$count = 76049;
	#10 counter$count = 76050;
	#10 counter$count = 76051;
	#10 counter$count = 76052;
	#10 counter$count = 76053;
	#10 counter$count = 76054;
	#10 counter$count = 76055;
	#10 counter$count = 76056;
	#10 counter$count = 76057;
	#10 counter$count = 76058;
	#10 counter$count = 76059;
	#10 counter$count = 76060;
	#10 counter$count = 76061;
	#10 counter$count = 76062;
	#10 counter$count = 76063;
	#10 counter$count = 76064;
	#10 counter$count = 76065;
	#10 counter$count = 76066;
	#10 counter$count = 76067;
	#10 counter$count = 76068;
	#10 counter$count = 76069;
	#10 counter$count = 76070;
	#10 counter$count = 76071;
	#10 counter$count = 76072;
	#10 counter$count = 76073;
	#10 counter$count = 76074;
	#10 counter$count = 76075;
	#10 counter$count = 76076;
	#10 counter$count = 76077;
	#10 counter$count = 76078;
	#10 counter$count = 76079;
	#10 counter$count = 76080;
	#10 counter$count = 76081;
	#10 counter$count = 76082;
	#10 counter$count = 76083;
	#10 counter$count = 76084;
	#10 counter$count = 76085;
	#10 counter$count = 76086;
	#10 counter$count = 76087;
	#10 counter$count = 76088;
	#10 counter$count = 76089;
	#10 counter$count = 76090;
	#10 counter$count = 76091;
	#10 counter$count = 76092;
	#10 counter$count = 76093;
	#10 counter$count = 76094;
	#10 counter$count = 76095;
	#10 counter$count = 76096;
	#10 counter$count = 76097;
	#10 counter$count = 76098;
	#10 counter$count = 76099;
	#10 counter$count = 76100;
	#10 counter$count = 76101;
	#10 counter$count = 76102;
	#10 counter$count = 76103;
	#10 counter$count = 76104;
	#10 counter$count = 76105;
	#10 counter$count = 76106;
	#10 counter$count = 76107;
	#10 counter$count = 76108;
	#10 counter$count = 76109;
	#10 counter$count = 76110;
	#10 counter$count = 76111;
	#10 counter$count = 76112;
	#10 counter$count = 76113;
	#10 counter$count = 76114;
	#10 counter$count = 76115;
	#10 counter$count = 76116;
	#10 counter$count = 76117;
	#10 counter$count = 76118;
	#10 counter$count = 76119;
	#10 counter$count = 76120;
	#10 counter$count = 76121;
	#10 counter$count = 76122;
	#10 counter$count = 76123;
	#10 counter$count = 76124;
	#10 counter$count = 76125;
	#10 counter$count = 76126;
	#10 counter$count = 76127;
	#10 counter$count = 76128;
	#10 counter$count = 76129;
	#10 counter$count = 76130;
	#10 counter$count = 76131;
	#10 counter$count = 76132;
	#10 counter$count = 76133;
	#10 counter$count = 76134;
	#10 counter$count = 76135;
	#10 counter$count = 76136;
	#10 counter$count = 76137;
	#10 counter$count = 76138;
	#10 counter$count = 76139;
	#10 counter$count = 76140;
	#10 counter$count = 76141;
	#10 counter$count = 76142;
	#10 counter$count = 76143;
	#10 counter$count = 76144;
	#10 counter$count = 76145;
	#10 counter$count = 76146;
	#10 counter$count = 76147;
	#10 counter$count = 76148;
	#10 counter$count = 76149;
	#10 counter$count = 76150;
	#10 counter$count = 76151;
	#10 counter$count = 76152;
	#10 counter$count = 76153;
	#10 counter$count = 76154;
	#10 counter$count = 76155;
	#10 counter$count = 76156;
	#10 counter$count = 76157;
	#10 counter$count = 76158;
	#10 counter$count = 76159;
	#10 counter$count = 76160;
	#10 counter$count = 76161;
	#10 counter$count = 76162;
	#10 counter$count = 76163;
	#10 counter$count = 76164;
	#10 counter$count = 76165;
	#10 counter$count = 76166;
	#10 counter$count = 76167;
	#10 counter$count = 76168;
	#10 counter$count = 76169;
	#10 counter$count = 76170;
	#10 counter$count = 76171;
	#10 counter$count = 76172;
	#10 counter$count = 76173;
	#10 counter$count = 76174;
	#10 counter$count = 76175;
	#10 counter$count = 76176;
	#10 counter$count = 76177;
	#10 counter$count = 76178;
	#10 counter$count = 76179;
	#10 counter$count = 76180;
	#10 counter$count = 76181;
	#10 counter$count = 76182;
	#10 counter$count = 76183;
	#10 counter$count = 76184;
	#10 counter$count = 76185;
	#10 counter$count = 76186;
	#10 counter$count = 76187;
	#10 counter$count = 76188;
	#10 counter$count = 76189;
	#10 counter$count = 76190;
	#10 counter$count = 76191;
	#10 counter$count = 76192;
	#10 counter$count = 76193;
	#10 counter$count = 76194;
	#10 counter$count = 76195;
	#10 counter$count = 76196;
	#10 counter$count = 76197;
	#10 counter$count = 76198;
	#10 counter$count = 76199;
	#10 counter$count = 76200;
	#10 counter$count = 76201;
	#10 counter$count = 76202;
	#10 counter$count = 76203;
	#10 counter$count = 76204;
	#10 counter$count = 76205;
	#10 counter$count = 76206;
	#10 counter$count = 76207;
	#10 counter$count = 76208;
	#10 counter$count = 76209;
	#10 counter$count = 76210;
	#10 counter$count = 76211;
	#10 counter$count = 76212;
	#10 counter$count = 76213;
	#10 counter$count = 76214;
	#10 counter$count = 76215;
	#10 counter$count = 76216;
	#10 counter$count = 76217;
	#10 counter$count = 76218;
	#10 counter$count = 76219;
	#10 counter$count = 76220;
	#10 counter$count = 76221;
	#10 counter$count = 76222;
	#10 counter$count = 76223;
	#10 counter$count = 76224;
	#10 counter$count = 76225;
	#10 counter$count = 76226;
	#10 counter$count = 76227;
	#10 counter$count = 76228;
	#10 counter$count = 76229;
	#10 counter$count = 76230;
	#10 counter$count = 76231;
	#10 counter$count = 76232;
	#10 counter$count = 76233;
	#10 counter$count = 76234;
	#10 counter$count = 76235;
	#10 counter$count = 76236;
	#10 counter$count = 76237;
	#10 counter$count = 76238;
	#10 counter$count = 76239;
	#10 counter$count = 76240;
	#10 counter$count = 76241;
	#10 counter$count = 76242;
	#10 counter$count = 76243;
	#10 counter$count = 76244;
	#10 counter$count = 76245;
	#10 counter$count = 76246;
	#10 counter$count = 76247;
	#10 counter$count = 76248;
	#10 counter$count = 76249;
	#10 counter$count = 76250;
	#10 counter$count = 76251;
	#10 counter$count = 76252;
	#10 counter$count = 76253;
	#10 counter$count = 76254;
	#10 counter$count = 76255;
	#10 counter$count = 76256;
	#10 counter$count = 76257;
	#10 counter$count = 76258;
	#10 counter$count = 76259;
	#10 counter$count = 76260;
	#10 counter$count = 76261;
	#10 counter$count = 76262;
	#10 counter$count = 76263;
	#10 counter$count = 76264;
	#10 counter$count = 76265;
	#10 counter$count = 76266;
	#10 counter$count = 76267;
	#10 counter$count = 76268;
	#10 counter$count = 76269;
	#10 counter$count = 76270;
	#10 counter$count = 76271;
	#10 counter$count = 76272;
	#10 counter$count = 76273;
	#10 counter$count = 76274;
	#10 counter$count = 76275;
	#10 counter$count = 76276;
	#10 counter$count = 76277;
	#10 counter$count = 76278;
	#10 counter$count = 76279;
	#10 counter$count = 76280;
	#10 counter$count = 76281;
	#10 counter$count = 76282;
	#10 counter$count = 76283;
	#10 counter$count = 76284;
	#10 counter$count = 76285;
	#10 counter$count = 76286;
	#10 counter$count = 76287;
	#10 counter$count = 76288;
	#10 counter$count = 76289;
	#10 counter$count = 76290;
	#10 counter$count = 76291;
	#10 counter$count = 76292;
	#10 counter$count = 76293;
	#10 counter$count = 76294;
	#10 counter$count = 76295;
	#10 counter$count = 76296;
	#10 counter$count = 76297;
	#10 counter$count = 76298;
	#10 counter$count = 76299;
	#10 counter$count = 76300;
	#10 counter$count = 76301;
	#10 counter$count = 76302;
	#10 counter$count = 76303;
	#10 counter$count = 76304;
	#10 counter$count = 76305;
	#10 counter$count = 76306;
	#10 counter$count = 76307;
	#10 counter$count = 76308;
	#10 counter$count = 76309;
	#10 counter$count = 76310;
	#10 counter$count = 76311;
	#10 counter$count = 76312;
	#10 counter$count = 76313;
	#10 counter$count = 76314;
	#10 counter$count = 76315;
	#10 counter$count = 76316;
	#10 counter$count = 76317;
	#10 counter$count = 76318;
	#10 counter$count = 76319;
	#10 counter$count = 76320;
	#10 counter$count = 76321;
	#10 counter$count = 76322;
	#10 counter$count = 76323;
	#10 counter$count = 76324;
	#10 counter$count = 76325;
	#10 counter$count = 76326;
	#10 counter$count = 76327;
	#10 counter$count = 76328;
	#10 counter$count = 76329;
	#10 counter$count = 76330;
	#10 counter$count = 76331;
	#10 counter$count = 76332;
	#10 counter$count = 76333;
	#10 counter$count = 76334;
	#10 counter$count = 76335;
	#10 counter$count = 76336;
	#10 counter$count = 76337;
	#10 counter$count = 76338;
	#10 counter$count = 76339;
	#10 counter$count = 76340;
	#10 counter$count = 76341;
	#10 counter$count = 76342;
	#10 counter$count = 76343;
	#10 counter$count = 76344;
	#10 counter$count = 76345;
	#10 counter$count = 76346;
	#10 counter$count = 76347;
	#10 counter$count = 76348;
	#10 counter$count = 76349;
	#10 counter$count = 76350;
	#10 counter$count = 76351;
	#10 counter$count = 76352;
	#10 counter$count = 76353;
	#10 counter$count = 76354;
	#10 counter$count = 76355;
	#10 counter$count = 76356;
	#10 counter$count = 76357;
	#10 counter$count = 76358;
	#10 counter$count = 76359;
	#10 counter$count = 76360;
	#10 counter$count = 76361;
	#10 counter$count = 76362;
	#10 counter$count = 76363;
	#10 counter$count = 76364;
	#10 counter$count = 76365;
	#10 counter$count = 76366;
	#10 counter$count = 76367;
	#10 counter$count = 76368;
	#10 counter$count = 76369;
	#10 counter$count = 76370;
	#10 counter$count = 76371;
	#10 counter$count = 76372;
	#10 counter$count = 76373;
	#10 counter$count = 76374;
	#10 counter$count = 76375;
	#10 counter$count = 76376;
	#10 counter$count = 76377;
	#10 counter$count = 76378;
	#10 counter$count = 76379;
	#10 counter$count = 76380;
	#10 counter$count = 76381;
	#10 counter$count = 76382;
	#10 counter$count = 76383;
	#10 counter$count = 76384;
	#10 counter$count = 76385;
	#10 counter$count = 76386;
	#10 counter$count = 76387;
	#10 counter$count = 76388;
	#10 counter$count = 76389;
	#10 counter$count = 76390;
	#10 counter$count = 76391;
	#10 counter$count = 76392;
	#10 counter$count = 76393;
	#10 counter$count = 76394;
	#10 counter$count = 76395;
	#10 counter$count = 76396;
	#10 counter$count = 76397;
	#10 counter$count = 76398;
	#10 counter$count = 76399;
	#10 counter$count = 76400;
	#10 counter$count = 76401;
	#10 counter$count = 76402;
	#10 counter$count = 76403;
	#10 counter$count = 76404;
	#10 counter$count = 76405;
	#10 counter$count = 76406;
	#10 counter$count = 76407;
	#10 counter$count = 76408;
	#10 counter$count = 76409;
	#10 counter$count = 76410;
	#10 counter$count = 76411;
	#10 counter$count = 76412;
	#10 counter$count = 76413;
	#10 counter$count = 76414;
	#10 counter$count = 76415;
	#10 counter$count = 76416;
	#10 counter$count = 76417;
	#10 counter$count = 76418;
	#10 counter$count = 76419;
	#10 counter$count = 76420;
	#10 counter$count = 76421;
	#10 counter$count = 76422;
	#10 counter$count = 76423;
	#10 counter$count = 76424;
	#10 counter$count = 76425;
	#10 counter$count = 76426;
	#10 counter$count = 76427;
	#10 counter$count = 76428;
	#10 counter$count = 76429;
	#10 counter$count = 76430;
	#10 counter$count = 76431;
	#10 counter$count = 76432;
	#10 counter$count = 76433;
	#10 counter$count = 76434;
	#10 counter$count = 76435;
	#10 counter$count = 76436;
	#10 counter$count = 76437;
	#10 counter$count = 76438;
	#10 counter$count = 76439;
	#10 counter$count = 76440;
	#10 counter$count = 76441;
	#10 counter$count = 76442;
	#10 counter$count = 76443;
	#10 counter$count = 76444;
	#10 counter$count = 76445;
	#10 counter$count = 76446;
	#10 counter$count = 76447;
	#10 counter$count = 76448;
	#10 counter$count = 76449;
	#10 counter$count = 76450;
	#10 counter$count = 76451;
	#10 counter$count = 76452;
	#10 counter$count = 76453;
	#10 counter$count = 76454;
	#10 counter$count = 76455;
	#10 counter$count = 76456;
	#10 counter$count = 76457;
	#10 counter$count = 76458;
	#10 counter$count = 76459;
	#10 counter$count = 76460;
	#10 counter$count = 76461;
	#10 counter$count = 76462;
	#10 counter$count = 76463;
	#10 counter$count = 76464;
	#10 counter$count = 76465;
	#10 counter$count = 76466;
	#10 counter$count = 76467;
	#10 counter$count = 76468;
	#10 counter$count = 76469;
	#10 counter$count = 76470;
	#10 counter$count = 76471;
	#10 counter$count = 76472;
	#10 counter$count = 76473;
	#10 counter$count = 76474;
	#10 counter$count = 76475;
	#10 counter$count = 76476;
	#10 counter$count = 76477;
	#10 counter$count = 76478;
	#10 counter$count = 76479;
	#10 counter$count = 76480;
	#10 counter$count = 76481;
	#10 counter$count = 76482;
	#10 counter$count = 76483;
	#10 counter$count = 76484;
	#10 counter$count = 76485;
	#10 counter$count = 76486;
	#10 counter$count = 76487;
	#10 counter$count = 76488;
	#10 counter$count = 76489;
	#10 counter$count = 76490;
	#10 counter$count = 76491;
	#10 counter$count = 76492;
	#10 counter$count = 76493;
	#10 counter$count = 76494;
	#10 counter$count = 76495;
	#10 counter$count = 76496;
	#10 counter$count = 76497;
	#10 counter$count = 76498;
	#10 counter$count = 76499;
	#10 counter$count = 76500;
	#10 counter$count = 76501;
	#10 counter$count = 76502;
	#10 counter$count = 76503;
	#10 counter$count = 76504;
	#10 counter$count = 76505;
	#10 counter$count = 76506;
	#10 counter$count = 76507;
	#10 counter$count = 76508;
	#10 counter$count = 76509;
	#10 counter$count = 76510;
	#10 counter$count = 76511;
	#10 counter$count = 76512;
	#10 counter$count = 76513;
	#10 counter$count = 76514;
	#10 counter$count = 76515;
	#10 counter$count = 76516;
	#10 counter$count = 76517;
	#10 counter$count = 76518;
	#10 counter$count = 76519;
	#10 counter$count = 76520;
	#10 counter$count = 76521;
	#10 counter$count = 76522;
	#10 counter$count = 76523;
	#10 counter$count = 76524;
	#10 counter$count = 76525;
	#10 counter$count = 76526;
	#10 counter$count = 76527;
	#10 counter$count = 76528;
	#10 counter$count = 76529;
	#10 counter$count = 76530;
	#10 counter$count = 76531;
	#10 counter$count = 76532;
	#10 counter$count = 76533;
	#10 counter$count = 76534;
	#10 counter$count = 76535;
	#10 counter$count = 76536;
	#10 counter$count = 76537;
	#10 counter$count = 76538;
	#10 counter$count = 76539;
	#10 counter$count = 76540;
	#10 counter$count = 76541;
	#10 counter$count = 76542;
	#10 counter$count = 76543;
	#10 counter$count = 76544;
	#10 counter$count = 76545;
	#10 counter$count = 76546;
	#10 counter$count = 76547;
	#10 counter$count = 76548;
	#10 counter$count = 76549;
	#10 counter$count = 76550;
	#10 counter$count = 76551;
	#10 counter$count = 76552;
	#10 counter$count = 76553;
	#10 counter$count = 76554;
	#10 counter$count = 76555;
	#10 counter$count = 76556;
	#10 counter$count = 76557;
	#10 counter$count = 76558;
	#10 counter$count = 76559;
	#10 counter$count = 76560;
	#10 counter$count = 76561;
	#10 counter$count = 76562;
	#10 counter$count = 76563;
	#10 counter$count = 76564;
	#10 counter$count = 76565;
	#10 counter$count = 76566;
	#10 counter$count = 76567;
	#10 counter$count = 76568;
	#10 counter$count = 76569;
	#10 counter$count = 76570;
	#10 counter$count = 76571;
	#10 counter$count = 76572;
	#10 counter$count = 76573;
	#10 counter$count = 76574;
	#10 counter$count = 76575;
	#10 counter$count = 76576;
	#10 counter$count = 76577;
	#10 counter$count = 76578;
	#10 counter$count = 76579;
	#10 counter$count = 76580;
	#10 counter$count = 76581;
	#10 counter$count = 76582;
	#10 counter$count = 76583;
	#10 counter$count = 76584;
	#10 counter$count = 76585;
	#10 counter$count = 76586;
	#10 counter$count = 76587;
	#10 counter$count = 76588;
	#10 counter$count = 76589;
	#10 counter$count = 76590;
	#10 counter$count = 76591;
	#10 counter$count = 76592;
	#10 counter$count = 76593;
	#10 counter$count = 76594;
	#10 counter$count = 76595;
	#10 counter$count = 76596;
	#10 counter$count = 76597;
	#10 counter$count = 76598;
	#10 counter$count = 76599;
	#10 counter$count = 76600;
	#10 counter$count = 76601;
	#10 counter$count = 76602;
	#10 counter$count = 76603;
	#10 counter$count = 76604;
	#10 counter$count = 76605;
	#10 counter$count = 76606;
	#10 counter$count = 76607;
	#10 counter$count = 76608;
	#10 counter$count = 76609;
	#10 counter$count = 76610;
	#10 counter$count = 76611;
	#10 counter$count = 76612;
	#10 counter$count = 76613;
	#10 counter$count = 76614;
	#10 counter$count = 76615;
	#10 counter$count = 76616;
	#10 counter$count = 76617;
	#10 counter$count = 76618;
	#10 counter$count = 76619;
	#10 counter$count = 76620;
	#10 counter$count = 76621;
	#10 counter$count = 76622;
	#10 counter$count = 76623;
	#10 counter$count = 76624;
	#10 counter$count = 76625;
	#10 counter$count = 76626;
	#10 counter$count = 76627;
	#10 counter$count = 76628;
	#10 counter$count = 76629;
	#10 counter$count = 76630;
	#10 counter$count = 76631;
	#10 counter$count = 76632;
	#10 counter$count = 76633;
	#10 counter$count = 76634;
	#10 counter$count = 76635;
	#10 counter$count = 76636;
	#10 counter$count = 76637;
	#10 counter$count = 76638;
	#10 counter$count = 76639;
	#10 counter$count = 76640;
	#10 counter$count = 76641;
	#10 counter$count = 76642;
	#10 counter$count = 76643;
	#10 counter$count = 76644;
	#10 counter$count = 76645;
	#10 counter$count = 76646;
	#10 counter$count = 76647;
	#10 counter$count = 76648;
	#10 counter$count = 76649;
	#10 counter$count = 76650;
	#10 counter$count = 76651;
	#10 counter$count = 76652;
	#10 counter$count = 76653;
	#10 counter$count = 76654;
	#10 counter$count = 76655;
	#10 counter$count = 76656;
	#10 counter$count = 76657;
	#10 counter$count = 76658;
	#10 counter$count = 76659;
	#10 counter$count = 76660;
	#10 counter$count = 76661;
	#10 counter$count = 76662;
	#10 counter$count = 76663;
	#10 counter$count = 76664;
	#10 counter$count = 76665;
	#10 counter$count = 76666;
	#10 counter$count = 76667;
	#10 counter$count = 76668;
	#10 counter$count = 76669;
	#10 counter$count = 76670;
	#10 counter$count = 76671;
	#10 counter$count = 76672;
	#10 counter$count = 76673;
	#10 counter$count = 76674;
	#10 counter$count = 76675;
	#10 counter$count = 76676;
	#10 counter$count = 76677;
	#10 counter$count = 76678;
	#10 counter$count = 76679;
	#10 counter$count = 76680;
	#10 counter$count = 76681;
	#10 counter$count = 76682;
	#10 counter$count = 76683;
	#10 counter$count = 76684;
	#10 counter$count = 76685;
	#10 counter$count = 76686;
	#10 counter$count = 76687;
	#10 counter$count = 76688;
	#10 counter$count = 76689;
	#10 counter$count = 76690;
	#10 counter$count = 76691;
	#10 counter$count = 76692;
	#10 counter$count = 76693;
	#10 counter$count = 76694;
	#10 counter$count = 76695;
	#10 counter$count = 76696;
	#10 counter$count = 76697;
	#10 counter$count = 76698;
	#10 counter$count = 76699;
	#10 counter$count = 76700;
	#10 counter$count = 76701;
	#10 counter$count = 76702;
	#10 counter$count = 76703;
	#10 counter$count = 76704;
	#10 counter$count = 76705;
	#10 counter$count = 76706;
	#10 counter$count = 76707;
	#10 counter$count = 76708;
	#10 counter$count = 76709;
	#10 counter$count = 76710;
	#10 counter$count = 76711;
	#10 counter$count = 76712;
	#10 counter$count = 76713;
	#10 counter$count = 76714;
	#10 counter$count = 76715;
	#10 counter$count = 76716;
	#10 counter$count = 76717;
	#10 counter$count = 76718;
	#10 counter$count = 76719;
	#10 counter$count = 76720;
	#10 counter$count = 76721;
	#10 counter$count = 76722;
	#10 counter$count = 76723;
	#10 counter$count = 76724;
	#10 counter$count = 76725;
	#10 counter$count = 76726;
	#10 counter$count = 76727;
	#10 counter$count = 76728;
	#10 counter$count = 76729;
	#10 counter$count = 76730;
	#10 counter$count = 76731;
	#10 counter$count = 76732;
	#10 counter$count = 76733;
	#10 counter$count = 76734;
	#10 counter$count = 76735;
	#10 counter$count = 76736;
	#10 counter$count = 76737;
	#10 counter$count = 76738;
	#10 counter$count = 76739;
	#10 counter$count = 76740;
	#10 counter$count = 76741;
	#10 counter$count = 76742;
	#10 counter$count = 76743;
	#10 counter$count = 76744;
	#10 counter$count = 76745;
	#10 counter$count = 76746;
	#10 counter$count = 76747;
	#10 counter$count = 76748;
	#10 counter$count = 76749;
	#10 counter$count = 76750;
	#10 counter$count = 76751;
	#10 counter$count = 76752;
	#10 counter$count = 76753;
	#10 counter$count = 76754;
	#10 counter$count = 76755;
	#10 counter$count = 76756;
	#10 counter$count = 76757;
	#10 counter$count = 76758;
	#10 counter$count = 76759;
	#10 counter$count = 76760;
	#10 counter$count = 76761;
	#10 counter$count = 76762;
	#10 counter$count = 76763;
	#10 counter$count = 76764;
	#10 counter$count = 76765;
	#10 counter$count = 76766;
	#10 counter$count = 76767;
	#10 counter$count = 76768;
	#10 counter$count = 76769;
	#10 counter$count = 76770;
	#10 counter$count = 76771;
	#10 counter$count = 76772;
	#10 counter$count = 76773;
	#10 counter$count = 76774;
	#10 counter$count = 76775;
	#10 counter$count = 76776;
	#10 counter$count = 76777;
	#10 counter$count = 76778;
	#10 counter$count = 76779;
	#10 counter$count = 76780;
	#10 counter$count = 76781;
	#10 counter$count = 76782;
	#10 counter$count = 76783;
	#10 counter$count = 76784;
	#10 counter$count = 76785;
	#10 counter$count = 76786;
	#10 counter$count = 76787;
	#10 counter$count = 76788;
	#10 counter$count = 76789;
	#10 counter$count = 76790;
	#10 counter$count = 76791;
	#10 counter$count = 76792;
	#10 counter$count = 76793;
	#10 counter$count = 76794;
	#10 counter$count = 76795;
	#10 counter$count = 76796;
	#10 counter$count = 76797;
	#10 counter$count = 76798;
	#10 counter$count = 76799;
	#10 counter$count = 76800;
	#10 counter$count = 76801;
	#10 counter$count = 76802;
	#10 counter$count = 76803;
	#10 counter$count = 76804;
	#10 counter$count = 76805;
	#10 counter$count = 76806;
	#10 counter$count = 76807;
	#10 counter$count = 76808;
	#10 counter$count = 76809;
	#10 counter$count = 76810;
	#10 counter$count = 76811;
	#10 counter$count = 76812;
	#10 counter$count = 76813;
	#10 counter$count = 76814;
	#10 counter$count = 76815;
	#10 counter$count = 76816;
	#10 counter$count = 76817;
	#10 counter$count = 76818;
	#10 counter$count = 76819;
	#10 counter$count = 76820;
	#10 counter$count = 76821;
	#10 counter$count = 76822;
	#10 counter$count = 76823;
	#10 counter$count = 76824;
	#10 counter$count = 76825;
	#10 counter$count = 76826;
	#10 counter$count = 76827;
	#10 counter$count = 76828;
	#10 counter$count = 76829;
	#10 counter$count = 76830;
	#10 counter$count = 76831;
	#10 counter$count = 76832;
	#10 counter$count = 76833;
	#10 counter$count = 76834;
	#10 counter$count = 76835;
	#10 counter$count = 76836;
	#10 counter$count = 76837;
	#10 counter$count = 76838;
	#10 counter$count = 76839;
	#10 counter$count = 76840;
	#10 counter$count = 76841;
	#10 counter$count = 76842;
	#10 counter$count = 76843;
	#10 counter$count = 76844;
	#10 counter$count = 76845;
	#10 counter$count = 76846;
	#10 counter$count = 76847;
	#10 counter$count = 76848;
	#10 counter$count = 76849;
	#10 counter$count = 76850;
	#10 counter$count = 76851;
	#10 counter$count = 76852;
	#10 counter$count = 76853;
	#10 counter$count = 76854;
	#10 counter$count = 76855;
	#10 counter$count = 76856;
	#10 counter$count = 76857;
	#10 counter$count = 76858;
	#10 counter$count = 76859;
	#10 counter$count = 76860;
	#10 counter$count = 76861;
	#10 counter$count = 76862;
	#10 counter$count = 76863;
	#10 counter$count = 76864;
	#10 counter$count = 76865;
	#10 counter$count = 76866;
	#10 counter$count = 76867;
	#10 counter$count = 76868;
	#10 counter$count = 76869;
	#10 counter$count = 76870;
	#10 counter$count = 76871;
	#10 counter$count = 76872;
	#10 counter$count = 76873;
	#10 counter$count = 76874;
	#10 counter$count = 76875;
	#10 counter$count = 76876;
	#10 counter$count = 76877;
	#10 counter$count = 76878;
	#10 counter$count = 76879;
	#10 counter$count = 76880;
	#10 counter$count = 76881;
	#10 counter$count = 76882;
	#10 counter$count = 76883;
	#10 counter$count = 76884;
	#10 counter$count = 76885;
	#10 counter$count = 76886;
	#10 counter$count = 76887;
	#10 counter$count = 76888;
	#10 counter$count = 76889;
	#10 counter$count = 76890;
	#10 counter$count = 76891;
	#10 counter$count = 76892;
	#10 counter$count = 76893;
	#10 counter$count = 76894;
	#10 counter$count = 76895;
	#10 counter$count = 76896;
	#10 counter$count = 76897;
	#10 counter$count = 76898;
	#10 counter$count = 76899;
	#10 counter$count = 76900;
	#10 counter$count = 76901;
	#10 counter$count = 76902;
	#10 counter$count = 76903;
	#10 counter$count = 76904;
	#10 counter$count = 76905;
	#10 counter$count = 76906;
	#10 counter$count = 76907;
	#10 counter$count = 76908;
	#10 counter$count = 76909;
	#10 counter$count = 76910;
	#10 counter$count = 76911;
	#10 counter$count = 76912;
	#10 counter$count = 76913;
	#10 counter$count = 76914;
	#10 counter$count = 76915;
	#10 counter$count = 76916;
	#10 counter$count = 76917;
	#10 counter$count = 76918;
	#10 counter$count = 76919;
	#10 counter$count = 76920;
	#10 counter$count = 76921;
	#10 counter$count = 76922;
	#10 counter$count = 76923;
	#10 counter$count = 76924;
	#10 counter$count = 76925;
	#10 counter$count = 76926;
	#10 counter$count = 76927;
	#10 counter$count = 76928;
	#10 counter$count = 76929;
	#10 counter$count = 76930;
	#10 counter$count = 76931;
	#10 counter$count = 76932;
	#10 counter$count = 76933;
	#10 counter$count = 76934;
	#10 counter$count = 76935;
	#10 counter$count = 76936;
	#10 counter$count = 76937;
	#10 counter$count = 76938;
	#10 counter$count = 76939;
	#10 counter$count = 76940;
	#10 counter$count = 76941;
	#10 counter$count = 76942;
	#10 counter$count = 76943;
	#10 counter$count = 76944;
	#10 counter$count = 76945;
	#10 counter$count = 76946;
	#10 counter$count = 76947;
	#10 counter$count = 76948;
	#10 counter$count = 76949;
	#10 counter$count = 76950;
	#10 counter$count = 76951;
	#10 counter$count = 76952;
	#10 counter$count = 76953;
	#10 counter$count = 76954;
	#10 counter$count = 76955;
	#10 counter$count = 76956;
	#10 counter$count = 76957;
	#10 counter$count = 76958;
	#10 counter$count = 76959;
	#10 counter$count = 76960;
	#10 counter$count = 76961;
	#10 counter$count = 76962;
	#10 counter$count = 76963;
	#10 counter$count = 76964;
	#10 counter$count = 76965;
	#10 counter$count = 76966;
	#10 counter$count = 76967;
	#10 counter$count = 76968;
	#10 counter$count = 76969;
	#10 counter$count = 76970;
	#10 counter$count = 76971;
	#10 counter$count = 76972;
	#10 counter$count = 76973;
	#10 counter$count = 76974;
	#10 counter$count = 76975;
	#10 counter$count = 76976;
	#10 counter$count = 76977;
	#10 counter$count = 76978;
	#10 counter$count = 76979;
	#10 counter$count = 76980;
	#10 counter$count = 76981;
	#10 counter$count = 76982;
	#10 counter$count = 76983;
	#10 counter$count = 76984;
	#10 counter$count = 76985;
	#10 counter$count = 76986;
	#10 counter$count = 76987;
	#10 counter$count = 76988;
	#10 counter$count = 76989;
	#10 counter$count = 76990;
	#10 counter$count = 76991;
	#10 counter$count = 76992;
	#10 counter$count = 76993;
	#10 counter$count = 76994;
	#10 counter$count = 76995;
	#10 counter$count = 76996;
	#10 counter$count = 76997;
	#10 counter$count = 76998;
	#10 counter$count = 76999;
	#10 counter$count = 77000;
	#10 counter$count = 77001;
	#10 counter$count = 77002;
	#10 counter$count = 77003;
	#10 counter$count = 77004;
	#10 counter$count = 77005;
	#10 counter$count = 77006;
	#10 counter$count = 77007;
	#10 counter$count = 77008;
	#10 counter$count = 77009;
	#10 counter$count = 77010;
	#10 counter$count = 77011;
	#10 counter$count = 77012;
	#10 counter$count = 77013;
	#10 counter$count = 77014;
	#10 counter$count = 77015;
	#10 counter$count = 77016;
	#10 counter$count = 77017;
	#10 counter$count = 77018;
	#10 counter$count = 77019;
	#10 counter$count = 77020;
	#10 counter$count = 77021;
	#10 counter$count = 77022;
	#10 counter$count = 77023;
	#10 counter$count = 77024;
	#10 counter$count = 77025;
	#10 counter$count = 77026;
	#10 counter$count = 77027;
	#10 counter$count = 77028;
	#10 counter$count = 77029;
	#10 counter$count = 77030;
	#10 counter$count = 77031;
	#10 counter$count = 77032;
	#10 counter$count = 77033;
	#10 counter$count = 77034;
	#10 counter$count = 77035;
	#10 counter$count = 77036;
	#10 counter$count = 77037;
	#10 counter$count = 77038;
	#10 counter$count = 77039;
	#10 counter$count = 77040;
	#10 counter$count = 77041;
	#10 counter$count = 77042;
	#10 counter$count = 77043;
	#10 counter$count = 77044;
	#10 counter$count = 77045;
	#10 counter$count = 77046;
	#10 counter$count = 77047;
	#10 counter$count = 77048;
	#10 counter$count = 77049;
	#10 counter$count = 77050;
	#10 counter$count = 77051;
	#10 counter$count = 77052;
	#10 counter$count = 77053;
	#10 counter$count = 77054;
	#10 counter$count = 77055;
	#10 counter$count = 77056;
	#10 counter$count = 77057;
	#10 counter$count = 77058;
	#10 counter$count = 77059;
	#10 counter$count = 77060;
	#10 counter$count = 77061;
	#10 counter$count = 77062;
	#10 counter$count = 77063;
	#10 counter$count = 77064;
	#10 counter$count = 77065;
	#10 counter$count = 77066;
	#10 counter$count = 77067;
	#10 counter$count = 77068;
	#10 counter$count = 77069;
	#10 counter$count = 77070;
	#10 counter$count = 77071;
	#10 counter$count = 77072;
	#10 counter$count = 77073;
	#10 counter$count = 77074;
	#10 counter$count = 77075;
	#10 counter$count = 77076;
	#10 counter$count = 77077;
	#10 counter$count = 77078;
	#10 counter$count = 77079;
	#10 counter$count = 77080;
	#10 counter$count = 77081;
	#10 counter$count = 77082;
	#10 counter$count = 77083;
	#10 counter$count = 77084;
	#10 counter$count = 77085;
	#10 counter$count = 77086;
	#10 counter$count = 77087;
	#10 counter$count = 77088;
	#10 counter$count = 77089;
	#10 counter$count = 77090;
	#10 counter$count = 77091;
	#10 counter$count = 77092;
	#10 counter$count = 77093;
	#10 counter$count = 77094;
	#10 counter$count = 77095;
	#10 counter$count = 77096;
	#10 counter$count = 77097;
	#10 counter$count = 77098;
	#10 counter$count = 77099;
	#10 counter$count = 77100;
	#10 counter$count = 77101;
	#10 counter$count = 77102;
	#10 counter$count = 77103;
	#10 counter$count = 77104;
	#10 counter$count = 77105;
	#10 counter$count = 77106;
	#10 counter$count = 77107;
	#10 counter$count = 77108;
	#10 counter$count = 77109;
	#10 counter$count = 77110;
	#10 counter$count = 77111;
	#10 counter$count = 77112;
	#10 counter$count = 77113;
	#10 counter$count = 77114;
	#10 counter$count = 77115;
	#10 counter$count = 77116;
	#10 counter$count = 77117;
	#10 counter$count = 77118;
	#10 counter$count = 77119;
	#10 counter$count = 77120;
	#10 counter$count = 77121;
	#10 counter$count = 77122;
	#10 counter$count = 77123;
	#10 counter$count = 77124;
	#10 counter$count = 77125;
	#10 counter$count = 77126;
	#10 counter$count = 77127;
	#10 counter$count = 77128;
	#10 counter$count = 77129;
	#10 counter$count = 77130;
	#10 counter$count = 77131;
	#10 counter$count = 77132;
	#10 counter$count = 77133;
	#10 counter$count = 77134;
	#10 counter$count = 77135;
	#10 counter$count = 77136;
	#10 counter$count = 77137;
	#10 counter$count = 77138;
	#10 counter$count = 77139;
	#10 counter$count = 77140;
	#10 counter$count = 77141;
	#10 counter$count = 77142;
	#10 counter$count = 77143;
	#10 counter$count = 77144;
	#10 counter$count = 77145;
	#10 counter$count = 77146;
	#10 counter$count = 77147;
	#10 counter$count = 77148;
	#10 counter$count = 77149;
	#10 counter$count = 77150;
	#10 counter$count = 77151;
	#10 counter$count = 77152;
	#10 counter$count = 77153;
	#10 counter$count = 77154;
	#10 counter$count = 77155;
	#10 counter$count = 77156;
	#10 counter$count = 77157;
	#10 counter$count = 77158;
	#10 counter$count = 77159;
	#10 counter$count = 77160;
	#10 counter$count = 77161;
	#10 counter$count = 77162;
	#10 counter$count = 77163;
	#10 counter$count = 77164;
	#10 counter$count = 77165;
	#10 counter$count = 77166;
	#10 counter$count = 77167;
	#10 counter$count = 77168;
	#10 counter$count = 77169;
	#10 counter$count = 77170;
	#10 counter$count = 77171;
	#10 counter$count = 77172;
	#10 counter$count = 77173;
	#10 counter$count = 77174;
	#10 counter$count = 77175;
	#10 counter$count = 77176;
	#10 counter$count = 77177;
	#10 counter$count = 77178;
	#10 counter$count = 77179;
	#10 counter$count = 77180;
	#10 counter$count = 77181;
	#10 counter$count = 77182;
	#10 counter$count = 77183;
	#10 counter$count = 77184;
	#10 counter$count = 77185;
	#10 counter$count = 77186;
	#10 counter$count = 77187;
	#10 counter$count = 77188;
	#10 counter$count = 77189;
	#10 counter$count = 77190;
	#10 counter$count = 77191;
	#10 counter$count = 77192;
	#10 counter$count = 77193;
	#10 counter$count = 77194;
	#10 counter$count = 77195;
	#10 counter$count = 77196;
	#10 counter$count = 77197;
	#10 counter$count = 77198;
	#10 counter$count = 77199;
	#10 counter$count = 77200;
	#10 counter$count = 77201;
	#10 counter$count = 77202;
	#10 counter$count = 77203;
	#10 counter$count = 77204;
	#10 counter$count = 77205;
	#10 counter$count = 77206;
	#10 counter$count = 77207;
	#10 counter$count = 77208;
	#10 counter$count = 77209;
	#10 counter$count = 77210;
	#10 counter$count = 77211;
	#10 counter$count = 77212;
	#10 counter$count = 77213;
	#10 counter$count = 77214;
	#10 counter$count = 77215;
	#10 counter$count = 77216;
	#10 counter$count = 77217;
	#10 counter$count = 77218;
	#10 counter$count = 77219;
	#10 counter$count = 77220;
	#10 counter$count = 77221;
	#10 counter$count = 77222;
	#10 counter$count = 77223;
	#10 counter$count = 77224;
	#10 counter$count = 77225;
	#10 counter$count = 77226;
	#10 counter$count = 77227;
	#10 counter$count = 77228;
	#10 counter$count = 77229;
	#10 counter$count = 77230;
	#10 counter$count = 77231;
	#10 counter$count = 77232;
	#10 counter$count = 77233;
	#10 counter$count = 77234;
	#10 counter$count = 77235;
	#10 counter$count = 77236;
	#10 counter$count = 77237;
	#10 counter$count = 77238;
	#10 counter$count = 77239;
	#10 counter$count = 77240;
	#10 counter$count = 77241;
	#10 counter$count = 77242;
	#10 counter$count = 77243;
	#10 counter$count = 77244;
	#10 counter$count = 77245;
	#10 counter$count = 77246;
	#10 counter$count = 77247;
	#10 counter$count = 77248;
	#10 counter$count = 77249;
	#10 counter$count = 77250;
	#10 counter$count = 77251;
	#10 counter$count = 77252;
	#10 counter$count = 77253;
	#10 counter$count = 77254;
	#10 counter$count = 77255;
	#10 counter$count = 77256;
	#10 counter$count = 77257;
	#10 counter$count = 77258;
	#10 counter$count = 77259;
	#10 counter$count = 77260;
	#10 counter$count = 77261;
	#10 counter$count = 77262;
	#10 counter$count = 77263;
	#10 counter$count = 77264;
	#10 counter$count = 77265;
	#10 counter$count = 77266;
	#10 counter$count = 77267;
	#10 counter$count = 77268;
	#10 counter$count = 77269;
	#10 counter$count = 77270;
	#10 counter$count = 77271;
	#10 counter$count = 77272;
	#10 counter$count = 77273;
	#10 counter$count = 77274;
	#10 counter$count = 77275;
	#10 counter$count = 77276;
	#10 counter$count = 77277;
	#10 counter$count = 77278;
	#10 counter$count = 77279;
	#10 counter$count = 77280;
	#10 counter$count = 77281;
	#10 counter$count = 77282;
	#10 counter$count = 77283;
	#10 counter$count = 77284;
	#10 counter$count = 77285;
	#10 counter$count = 77286;
	#10 counter$count = 77287;
	#10 counter$count = 77288;
	#10 counter$count = 77289;
	#10 counter$count = 77290;
	#10 counter$count = 77291;
	#10 counter$count = 77292;
	#10 counter$count = 77293;
	#10 counter$count = 77294;
	#10 counter$count = 77295;
	#10 counter$count = 77296;
	#10 counter$count = 77297;
	#10 counter$count = 77298;
	#10 counter$count = 77299;
	#10 counter$count = 77300;
	#10 counter$count = 77301;
	#10 counter$count = 77302;
	#10 counter$count = 77303;
	#10 counter$count = 77304;
	#10 counter$count = 77305;
	#10 counter$count = 77306;
	#10 counter$count = 77307;
	#10 counter$count = 77308;
	#10 counter$count = 77309;
	#10 counter$count = 77310;
	#10 counter$count = 77311;
	#10 counter$count = 77312;
	#10 counter$count = 77313;
	#10 counter$count = 77314;
	#10 counter$count = 77315;
	#10 counter$count = 77316;
	#10 counter$count = 77317;
	#10 counter$count = 77318;
	#10 counter$count = 77319;
	#10 counter$count = 77320;
	#10 counter$count = 77321;
	#10 counter$count = 77322;
	#10 counter$count = 77323;
	#10 counter$count = 77324;
	#10 counter$count = 77325;
	#10 counter$count = 77326;
	#10 counter$count = 77327;
	#10 counter$count = 77328;
	#10 counter$count = 77329;
	#10 counter$count = 77330;
	#10 counter$count = 77331;
	#10 counter$count = 77332;
	#10 counter$count = 77333;
	#10 counter$count = 77334;
	#10 counter$count = 77335;
	#10 counter$count = 77336;
	#10 counter$count = 77337;
	#10 counter$count = 77338;
	#10 counter$count = 77339;
	#10 counter$count = 77340;
	#10 counter$count = 77341;
	#10 counter$count = 77342;
	#10 counter$count = 77343;
	#10 counter$count = 77344;
	#10 counter$count = 77345;
	#10 counter$count = 77346;
	#10 counter$count = 77347;
	#10 counter$count = 77348;
	#10 counter$count = 77349;
	#10 counter$count = 77350;
	#10 counter$count = 77351;
	#10 counter$count = 77352;
	#10 counter$count = 77353;
	#10 counter$count = 77354;
	#10 counter$count = 77355;
	#10 counter$count = 77356;
	#10 counter$count = 77357;
	#10 counter$count = 77358;
	#10 counter$count = 77359;
	#10 counter$count = 77360;
	#10 counter$count = 77361;
	#10 counter$count = 77362;
	#10 counter$count = 77363;
	#10 counter$count = 77364;
	#10 counter$count = 77365;
	#10 counter$count = 77366;
	#10 counter$count = 77367;
	#10 counter$count = 77368;
	#10 counter$count = 77369;
	#10 counter$count = 77370;
	#10 counter$count = 77371;
	#10 counter$count = 77372;
	#10 counter$count = 77373;
	#10 counter$count = 77374;
	#10 counter$count = 77375;
	#10 counter$count = 77376;
	#10 counter$count = 77377;
	#10 counter$count = 77378;
	#10 counter$count = 77379;
	#10 counter$count = 77380;
	#10 counter$count = 77381;
	#10 counter$count = 77382;
	#10 counter$count = 77383;
	#10 counter$count = 77384;
	#10 counter$count = 77385;
	#10 counter$count = 77386;
	#10 counter$count = 77387;
	#10 counter$count = 77388;
	#10 counter$count = 77389;
	#10 counter$count = 77390;
	#10 counter$count = 77391;
	#10 counter$count = 77392;
	#10 counter$count = 77393;
	#10 counter$count = 77394;
	#10 counter$count = 77395;
	#10 counter$count = 77396;
	#10 counter$count = 77397;
	#10 counter$count = 77398;
	#10 counter$count = 77399;
	#10 counter$count = 77400;
	#10 counter$count = 77401;
	#10 counter$count = 77402;
	#10 counter$count = 77403;
	#10 counter$count = 77404;
	#10 counter$count = 77405;
	#10 counter$count = 77406;
	#10 counter$count = 77407;
	#10 counter$count = 77408;
	#10 counter$count = 77409;
	#10 counter$count = 77410;
	#10 counter$count = 77411;
	#10 counter$count = 77412;
	#10 counter$count = 77413;
	#10 counter$count = 77414;
	#10 counter$count = 77415;
	#10 counter$count = 77416;
	#10 counter$count = 77417;
	#10 counter$count = 77418;
	#10 counter$count = 77419;
	#10 counter$count = 77420;
	#10 counter$count = 77421;
	#10 counter$count = 77422;
	#10 counter$count = 77423;
	#10 counter$count = 77424;
	#10 counter$count = 77425;
	#10 counter$count = 77426;
	#10 counter$count = 77427;
	#10 counter$count = 77428;
	#10 counter$count = 77429;
	#10 counter$count = 77430;
	#10 counter$count = 77431;
	#10 counter$count = 77432;
	#10 counter$count = 77433;
	#10 counter$count = 77434;
	#10 counter$count = 77435;
	#10 counter$count = 77436;
	#10 counter$count = 77437;
	#10 counter$count = 77438;
	#10 counter$count = 77439;
	#10 counter$count = 77440;
	#10 counter$count = 77441;
	#10 counter$count = 77442;
	#10 counter$count = 77443;
	#10 counter$count = 77444;
	#10 counter$count = 77445;
	#10 counter$count = 77446;
	#10 counter$count = 77447;
	#10 counter$count = 77448;
	#10 counter$count = 77449;
	#10 counter$count = 77450;
	#10 counter$count = 77451;
	#10 counter$count = 77452;
	#10 counter$count = 77453;
	#10 counter$count = 77454;
	#10 counter$count = 77455;
	#10 counter$count = 77456;
	#10 counter$count = 77457;
	#10 counter$count = 77458;
	#10 counter$count = 77459;
	#10 counter$count = 77460;
	#10 counter$count = 77461;
	#10 counter$count = 77462;
	#10 counter$count = 77463;
	#10 counter$count = 77464;
	#10 counter$count = 77465;
	#10 counter$count = 77466;
	#10 counter$count = 77467;
	#10 counter$count = 77468;
	#10 counter$count = 77469;
	#10 counter$count = 77470;
	#10 counter$count = 77471;
	#10 counter$count = 77472;
	#10 counter$count = 77473;
	#10 counter$count = 77474;
	#10 counter$count = 77475;
	#10 counter$count = 77476;
	#10 counter$count = 77477;
	#10 counter$count = 77478;
	#10 counter$count = 77479;
	#10 counter$count = 77480;
	#10 counter$count = 77481;
	#10 counter$count = 77482;
	#10 counter$count = 77483;
	#10 counter$count = 77484;
	#10 counter$count = 77485;
	#10 counter$count = 77486;
	#10 counter$count = 77487;
	#10 counter$count = 77488;
	#10 counter$count = 77489;
	#10 counter$count = 77490;
	#10 counter$count = 77491;
	#10 counter$count = 77492;
	#10 counter$count = 77493;
	#10 counter$count = 77494;
	#10 counter$count = 77495;
	#10 counter$count = 77496;
	#10 counter$count = 77497;
	#10 counter$count = 77498;
	#10 counter$count = 77499;
	#10 counter$count = 77500;
	#10 counter$count = 77501;
	#10 counter$count = 77502;
	#10 counter$count = 77503;
	#10 counter$count = 77504;
	#10 counter$count = 77505;
	#10 counter$count = 77506;
	#10 counter$count = 77507;
	#10 counter$count = 77508;
	#10 counter$count = 77509;
	#10 counter$count = 77510;
	#10 counter$count = 77511;
	#10 counter$count = 77512;
	#10 counter$count = 77513;
	#10 counter$count = 77514;
	#10 counter$count = 77515;
	#10 counter$count = 77516;
	#10 counter$count = 77517;
	#10 counter$count = 77518;
	#10 counter$count = 77519;
	#10 counter$count = 77520;
	#10 counter$count = 77521;
	#10 counter$count = 77522;
	#10 counter$count = 77523;
	#10 counter$count = 77524;
	#10 counter$count = 77525;
	#10 counter$count = 77526;
	#10 counter$count = 77527;
	#10 counter$count = 77528;
	#10 counter$count = 77529;
	#10 counter$count = 77530;
	#10 counter$count = 77531;
	#10 counter$count = 77532;
	#10 counter$count = 77533;
	#10 counter$count = 77534;
	#10 counter$count = 77535;
	#10 counter$count = 77536;
	#10 counter$count = 77537;
	#10 counter$count = 77538;
	#10 counter$count = 77539;
	#10 counter$count = 77540;
	#10 counter$count = 77541;
	#10 counter$count = 77542;
	#10 counter$count = 77543;
	#10 counter$count = 77544;
	#10 counter$count = 77545;
	#10 counter$count = 77546;
	#10 counter$count = 77547;
	#10 counter$count = 77548;
	#10 counter$count = 77549;
	#10 counter$count = 77550;
	#10 counter$count = 77551;
	#10 counter$count = 77552;
	#10 counter$count = 77553;
	#10 counter$count = 77554;
	#10 counter$count = 77555;
	#10 counter$count = 77556;
	#10 counter$count = 77557;
	#10 counter$count = 77558;
	#10 counter$count = 77559;
	#10 counter$count = 77560;
	#10 counter$count = 77561;
	#10 counter$count = 77562;
	#10 counter$count = 77563;
	#10 counter$count = 77564;
	#10 counter$count = 77565;
	#10 counter$count = 77566;
	#10 counter$count = 77567;
	#10 counter$count = 77568;
	#10 counter$count = 77569;
	#10 counter$count = 77570;
	#10 counter$count = 77571;
	#10 counter$count = 77572;
	#10 counter$count = 77573;
	#10 counter$count = 77574;
	#10 counter$count = 77575;
	#10 counter$count = 77576;
	#10 counter$count = 77577;
	#10 counter$count = 77578;
	#10 counter$count = 77579;
	#10 counter$count = 77580;
	#10 counter$count = 77581;
	#10 counter$count = 77582;
	#10 counter$count = 77583;
	#10 counter$count = 77584;
	#10 counter$count = 77585;
	#10 counter$count = 77586;
	#10 counter$count = 77587;
	#10 counter$count = 77588;
	#10 counter$count = 77589;
	#10 counter$count = 77590;
	#10 counter$count = 77591;
	#10 counter$count = 77592;
	#10 counter$count = 77593;
	#10 counter$count = 77594;
	#10 counter$count = 77595;
	#10 counter$count = 77596;
	#10 counter$count = 77597;
	#10 counter$count = 77598;
	#10 counter$count = 77599;
	#10 counter$count = 77600;
	#10 counter$count = 77601;
	#10 counter$count = 77602;
	#10 counter$count = 77603;
	#10 counter$count = 77604;
	#10 counter$count = 77605;
	#10 counter$count = 77606;
	#10 counter$count = 77607;
	#10 counter$count = 77608;
	#10 counter$count = 77609;
	#10 counter$count = 77610;
	#10 counter$count = 77611;
	#10 counter$count = 77612;
	#10 counter$count = 77613;
	#10 counter$count = 77614;
	#10 counter$count = 77615;
	#10 counter$count = 77616;
	#10 counter$count = 77617;
	#10 counter$count = 77618;
	#10 counter$count = 77619;
	#10 counter$count = 77620;
	#10 counter$count = 77621;
	#10 counter$count = 77622;
	#10 counter$count = 77623;
	#10 counter$count = 77624;
	#10 counter$count = 77625;
	#10 counter$count = 77626;
	#10 counter$count = 77627;
	#10 counter$count = 77628;
	#10 counter$count = 77629;
	#10 counter$count = 77630;
	#10 counter$count = 77631;
	#10 counter$count = 77632;
	#10 counter$count = 77633;
	#10 counter$count = 77634;
	#10 counter$count = 77635;
	#10 counter$count = 77636;
	#10 counter$count = 77637;
	#10 counter$count = 77638;
	#10 counter$count = 77639;
	#10 counter$count = 77640;
	#10 counter$count = 77641;
	#10 counter$count = 77642;
	#10 counter$count = 77643;
	#10 counter$count = 77644;
	#10 counter$count = 77645;
	#10 counter$count = 77646;
	#10 counter$count = 77647;
	#10 counter$count = 77648;
	#10 counter$count = 77649;
	#10 counter$count = 77650;
	#10 counter$count = 77651;
	#10 counter$count = 77652;
	#10 counter$count = 77653;
	#10 counter$count = 77654;
	#10 counter$count = 77655;
	#10 counter$count = 77656;
	#10 counter$count = 77657;
	#10 counter$count = 77658;
	#10 counter$count = 77659;
	#10 counter$count = 77660;
	#10 counter$count = 77661;
	#10 counter$count = 77662;
	#10 counter$count = 77663;
	#10 counter$count = 77664;
	#10 counter$count = 77665;
	#10 counter$count = 77666;
	#10 counter$count = 77667;
	#10 counter$count = 77668;
	#10 counter$count = 77669;
	#10 counter$count = 77670;
	#10 counter$count = 77671;
	#10 counter$count = 77672;
	#10 counter$count = 77673;
	#10 counter$count = 77674;
	#10 counter$count = 77675;
	#10 counter$count = 77676;
	#10 counter$count = 77677;
	#10 counter$count = 77678;
	#10 counter$count = 77679;
	#10 counter$count = 77680;
	#10 counter$count = 77681;
	#10 counter$count = 77682;
	#10 counter$count = 77683;
	#10 counter$count = 77684;
	#10 counter$count = 77685;
	#10 counter$count = 77686;
	#10 counter$count = 77687;
	#10 counter$count = 77688;
	#10 counter$count = 77689;
	#10 counter$count = 77690;
	#10 counter$count = 77691;
	#10 counter$count = 77692;
	#10 counter$count = 77693;
	#10 counter$count = 77694;
	#10 counter$count = 77695;
	#10 counter$count = 77696;
	#10 counter$count = 77697;
	#10 counter$count = 77698;
	#10 counter$count = 77699;
	#10 counter$count = 77700;
	#10 counter$count = 77701;
	#10 counter$count = 77702;
	#10 counter$count = 77703;
	#10 counter$count = 77704;
	#10 counter$count = 77705;
	#10 counter$count = 77706;
	#10 counter$count = 77707;
	#10 counter$count = 77708;
	#10 counter$count = 77709;
	#10 counter$count = 77710;
	#10 counter$count = 77711;
	#10 counter$count = 77712;
	#10 counter$count = 77713;
	#10 counter$count = 77714;
	#10 counter$count = 77715;
	#10 counter$count = 77716;
	#10 counter$count = 77717;
	#10 counter$count = 77718;
	#10 counter$count = 77719;
	#10 counter$count = 77720;
	#10 counter$count = 77721;
	#10 counter$count = 77722;
	#10 counter$count = 77723;
	#10 counter$count = 77724;
	#10 counter$count = 77725;
	#10 counter$count = 77726;
	#10 counter$count = 77727;
	#10 counter$count = 77728;
	#10 counter$count = 77729;
	#10 counter$count = 77730;
	#10 counter$count = 77731;
	#10 counter$count = 77732;
	#10 counter$count = 77733;
	#10 counter$count = 77734;
	#10 counter$count = 77735;
	#10 counter$count = 77736;
	#10 counter$count = 77737;
	#10 counter$count = 77738;
	#10 counter$count = 77739;
	#10 counter$count = 77740;
	#10 counter$count = 77741;
	#10 counter$count = 77742;
	#10 counter$count = 77743;
	#10 counter$count = 77744;
	#10 counter$count = 77745;
	#10 counter$count = 77746;
	#10 counter$count = 77747;
	#10 counter$count = 77748;
	#10 counter$count = 77749;
	#10 counter$count = 77750;
	#10 counter$count = 77751;
	#10 counter$count = 77752;
	#10 counter$count = 77753;
	#10 counter$count = 77754;
	#10 counter$count = 77755;
	#10 counter$count = 77756;
	#10 counter$count = 77757;
	#10 counter$count = 77758;
	#10 counter$count = 77759;
	#10 counter$count = 77760;
	#10 counter$count = 77761;
	#10 counter$count = 77762;
	#10 counter$count = 77763;
	#10 counter$count = 77764;
	#10 counter$count = 77765;
	#10 counter$count = 77766;
	#10 counter$count = 77767;
	#10 counter$count = 77768;
	#10 counter$count = 77769;
	#10 counter$count = 77770;
	#10 counter$count = 77771;
	#10 counter$count = 77772;
	#10 counter$count = 77773;
	#10 counter$count = 77774;
	#10 counter$count = 77775;
	#10 counter$count = 77776;
	#10 counter$count = 77777;
	#10 counter$count = 77778;
	#10 counter$count = 77779;
	#10 counter$count = 77780;
	#10 counter$count = 77781;
	#10 counter$count = 77782;
	#10 counter$count = 77783;
	#10 counter$count = 77784;
	#10 counter$count = 77785;
	#10 counter$count = 77786;
	#10 counter$count = 77787;
	#10 counter$count = 77788;
	#10 counter$count = 77789;
	#10 counter$count = 77790;
	#10 counter$count = 77791;
	#10 counter$count = 77792;
	#10 counter$count = 77793;
	#10 counter$count = 77794;
	#10 counter$count = 77795;
	#10 counter$count = 77796;
	#10 counter$count = 77797;
	#10 counter$count = 77798;
	#10 counter$count = 77799;
	#10 counter$count = 77800;
	#10 counter$count = 77801;
	#10 counter$count = 77802;
	#10 counter$count = 77803;
	#10 counter$count = 77804;
	#10 counter$count = 77805;
	#10 counter$count = 77806;
	#10 counter$count = 77807;
	#10 counter$count = 77808;
	#10 counter$count = 77809;
	#10 counter$count = 77810;
	#10 counter$count = 77811;
	#10 counter$count = 77812;
	#10 counter$count = 77813;
	#10 counter$count = 77814;
	#10 counter$count = 77815;
	#10 counter$count = 77816;
	#10 counter$count = 77817;
	#10 counter$count = 77818;
	#10 counter$count = 77819;
	#10 counter$count = 77820;
	#10 counter$count = 77821;
	#10 counter$count = 77822;
	#10 counter$count = 77823;
	#10 counter$count = 77824;
	#10 counter$count = 77825;
	#10 counter$count = 77826;
	#10 counter$count = 77827;
	#10 counter$count = 77828;
	#10 counter$count = 77829;
	#10 counter$count = 77830;
	#10 counter$count = 77831;
	#10 counter$count = 77832;
	#10 counter$count = 77833;
	#10 counter$count = 77834;
	#10 counter$count = 77835;
	#10 counter$count = 77836;
	#10 counter$count = 77837;
	#10 counter$count = 77838;
	#10 counter$count = 77839;
	#10 counter$count = 77840;
	#10 counter$count = 77841;
	#10 counter$count = 77842;
	#10 counter$count = 77843;
	#10 counter$count = 77844;
	#10 counter$count = 77845;
	#10 counter$count = 77846;
	#10 counter$count = 77847;
	#10 counter$count = 77848;
	#10 counter$count = 77849;
	#10 counter$count = 77850;
	#10 counter$count = 77851;
	#10 counter$count = 77852;
	#10 counter$count = 77853;
	#10 counter$count = 77854;
	#10 counter$count = 77855;
	#10 counter$count = 77856;
	#10 counter$count = 77857;
	#10 counter$count = 77858;
	#10 counter$count = 77859;
	#10 counter$count = 77860;
	#10 counter$count = 77861;
	#10 counter$count = 77862;
	#10 counter$count = 77863;
	#10 counter$count = 77864;
	#10 counter$count = 77865;
	#10 counter$count = 77866;
	#10 counter$count = 77867;
	#10 counter$count = 77868;
	#10 counter$count = 77869;
	#10 counter$count = 77870;
	#10 counter$count = 77871;
	#10 counter$count = 77872;
	#10 counter$count = 77873;
	#10 counter$count = 77874;
	#10 counter$count = 77875;
	#10 counter$count = 77876;
	#10 counter$count = 77877;
	#10 counter$count = 77878;
	#10 counter$count = 77879;
	#10 counter$count = 77880;
	#10 counter$count = 77881;
	#10 counter$count = 77882;
	#10 counter$count = 77883;
	#10 counter$count = 77884;
	#10 counter$count = 77885;
	#10 counter$count = 77886;
	#10 counter$count = 77887;
	#10 counter$count = 77888;
	#10 counter$count = 77889;
	#10 counter$count = 77890;
	#10 counter$count = 77891;
	#10 counter$count = 77892;
	#10 counter$count = 77893;
	#10 counter$count = 77894;
	#10 counter$count = 77895;
	#10 counter$count = 77896;
	#10 counter$count = 77897;
	#10 counter$count = 77898;
	#10 counter$count = 77899;
	#10 counter$count = 77900;
	#10 counter$count = 77901;
	#10 counter$count = 77902;
	#10 counter$count = 77903;
	#10 counter$count = 77904;
	#10 counter$count = 77905;
	#10 counter$count = 77906;
	#10 counter$count = 77907;
	#10 counter$count = 77908;
	#10 counter$count = 77909;
	#10 counter$count = 77910;
	#10 counter$count = 77911;
	#10 counter$count = 77912;
	#10 counter$count = 77913;
	#10 counter$count = 77914;
	#10 counter$count = 77915;
	#10 counter$count = 77916;
	#10 counter$count = 77917;
	#10 counter$count = 77918;
	#10 counter$count = 77919;
	#10 counter$count = 77920;
	#10 counter$count = 77921;
	#10 counter$count = 77922;
	#10 counter$count = 77923;
	#10 counter$count = 77924;
	#10 counter$count = 77925;
	#10 counter$count = 77926;
	#10 counter$count = 77927;
	#10 counter$count = 77928;
	#10 counter$count = 77929;
	#10 counter$count = 77930;
	#10 counter$count = 77931;
	#10 counter$count = 77932;
	#10 counter$count = 77933;
	#10 counter$count = 77934;
	#10 counter$count = 77935;
	#10 counter$count = 77936;
	#10 counter$count = 77937;
	#10 counter$count = 77938;
	#10 counter$count = 77939;
	#10 counter$count = 77940;
	#10 counter$count = 77941;
	#10 counter$count = 77942;
	#10 counter$count = 77943;
	#10 counter$count = 77944;
	#10 counter$count = 77945;
	#10 counter$count = 77946;
	#10 counter$count = 77947;
	#10 counter$count = 77948;
	#10 counter$count = 77949;
	#10 counter$count = 77950;
	#10 counter$count = 77951;
	#10 counter$count = 77952;
	#10 counter$count = 77953;
	#10 counter$count = 77954;
	#10 counter$count = 77955;
	#10 counter$count = 77956;
	#10 counter$count = 77957;
	#10 counter$count = 77958;
	#10 counter$count = 77959;
	#10 counter$count = 77960;
	#10 counter$count = 77961;
	#10 counter$count = 77962;
	#10 counter$count = 77963;
	#10 counter$count = 77964;
	#10 counter$count = 77965;
	#10 counter$count = 77966;
	#10 counter$count = 77967;
	#10 counter$count = 77968;
	#10 counter$count = 77969;
	#10 counter$count = 77970;
	#10 counter$count = 77971;
	#10 counter$count = 77972;
	#10 counter$count = 77973;
	#10 counter$count = 77974;
	#10 counter$count = 77975;
	#10 counter$count = 77976;
	#10 counter$count = 77977;
	#10 counter$count = 77978;
	#10 counter$count = 77979;
	#10 counter$count = 77980;
	#10 counter$count = 77981;
	#10 counter$count = 77982;
	#10 counter$count = 77983;
	#10 counter$count = 77984;
	#10 counter$count = 77985;
	#10 counter$count = 77986;
	#10 counter$count = 77987;
	#10 counter$count = 77988;
	#10 counter$count = 77989;
	#10 counter$count = 77990;
	#10 counter$count = 77991;
	#10 counter$count = 77992;
	#10 counter$count = 77993;
	#10 counter$count = 77994;
	#10 counter$count = 77995;
	#10 counter$count = 77996;
	#10 counter$count = 77997;
	#10 counter$count = 77998;
	#10 counter$count = 77999;
	#10 counter$count = 78000;
	#10 counter$count = 78001;
	#10 counter$count = 78002;
	#10 counter$count = 78003;
	#10 counter$count = 78004;
	#10 counter$count = 78005;
	#10 counter$count = 78006;
	#10 counter$count = 78007;
	#10 counter$count = 78008;
	#10 counter$count = 78009;
	#10 counter$count = 78010;
	#10 counter$count = 78011;
	#10 counter$count = 78012;
	#10 counter$count = 78013;
	#10 counter$count = 78014;
	#10 counter$count = 78015;
	#10 counter$count = 78016;
	#10 counter$count = 78017;
	#10 counter$count = 78018;
	#10 counter$count = 78019;
	#10 counter$count = 78020;
	#10 counter$count = 78021;
	#10 counter$count = 78022;
	#10 counter$count = 78023;
	#10 counter$count = 78024;
	#10 counter$count = 78025;
	#10 counter$count = 78026;
	#10 counter$count = 78027;
	#10 counter$count = 78028;
	#10 counter$count = 78029;
	#10 counter$count = 78030;
	#10 counter$count = 78031;
	#10 counter$count = 78032;
	#10 counter$count = 78033;
	#10 counter$count = 78034;
	#10 counter$count = 78035;
	#10 counter$count = 78036;
	#10 counter$count = 78037;
	#10 counter$count = 78038;
	#10 counter$count = 78039;
	#10 counter$count = 78040;
	#10 counter$count = 78041;
	#10 counter$count = 78042;
	#10 counter$count = 78043;
	#10 counter$count = 78044;
	#10 counter$count = 78045;
	#10 counter$count = 78046;
	#10 counter$count = 78047;
	#10 counter$count = 78048;
	#10 counter$count = 78049;
	#10 counter$count = 78050;
	#10 counter$count = 78051;
	#10 counter$count = 78052;
	#10 counter$count = 78053;
	#10 counter$count = 78054;
	#10 counter$count = 78055;
	#10 counter$count = 78056;
	#10 counter$count = 78057;
	#10 counter$count = 78058;
	#10 counter$count = 78059;
	#10 counter$count = 78060;
	#10 counter$count = 78061;
	#10 counter$count = 78062;
	#10 counter$count = 78063;
	#10 counter$count = 78064;
	#10 counter$count = 78065;
	#10 counter$count = 78066;
	#10 counter$count = 78067;
	#10 counter$count = 78068;
	#10 counter$count = 78069;
	#10 counter$count = 78070;
	#10 counter$count = 78071;
	#10 counter$count = 78072;
	#10 counter$count = 78073;
	#10 counter$count = 78074;
	#10 counter$count = 78075;
	#10 counter$count = 78076;
	#10 counter$count = 78077;
	#10 counter$count = 78078;
	#10 counter$count = 78079;
	#10 counter$count = 78080;
	#10 counter$count = 78081;
	#10 counter$count = 78082;
	#10 counter$count = 78083;
	#10 counter$count = 78084;
	#10 counter$count = 78085;
	#10 counter$count = 78086;
	#10 counter$count = 78087;
	#10 counter$count = 78088;
	#10 counter$count = 78089;
	#10 counter$count = 78090;
	#10 counter$count = 78091;
	#10 counter$count = 78092;
	#10 counter$count = 78093;
	#10 counter$count = 78094;
	#10 counter$count = 78095;
	#10 counter$count = 78096;
	#10 counter$count = 78097;
	#10 counter$count = 78098;
	#10 counter$count = 78099;
	#10 counter$count = 78100;
	#10 counter$count = 78101;
	#10 counter$count = 78102;
	#10 counter$count = 78103;
	#10 counter$count = 78104;
	#10 counter$count = 78105;
	#10 counter$count = 78106;
	#10 counter$count = 78107;
	#10 counter$count = 78108;
	#10 counter$count = 78109;
	#10 counter$count = 78110;
	#10 counter$count = 78111;
	#10 counter$count = 78112;
	#10 counter$count = 78113;
	#10 counter$count = 78114;
	#10 counter$count = 78115;
	#10 counter$count = 78116;
	#10 counter$count = 78117;
	#10 counter$count = 78118;
	#10 counter$count = 78119;
	#10 counter$count = 78120;
	#10 counter$count = 78121;
	#10 counter$count = 78122;
	#10 counter$count = 78123;
	#10 counter$count = 78124;
	#10 counter$count = 78125;
	#10 counter$count = 78126;
	#10 counter$count = 78127;
	#10 counter$count = 78128;
	#10 counter$count = 78129;
	#10 counter$count = 78130;
	#10 counter$count = 78131;
	#10 counter$count = 78132;
	#10 counter$count = 78133;
	#10 counter$count = 78134;
	#10 counter$count = 78135;
	#10 counter$count = 78136;
	#10 counter$count = 78137;
	#10 counter$count = 78138;
	#10 counter$count = 78139;
	#10 counter$count = 78140;
	#10 counter$count = 78141;
	#10 counter$count = 78142;
	#10 counter$count = 78143;
	#10 counter$count = 78144;
	#10 counter$count = 78145;
	#10 counter$count = 78146;
	#10 counter$count = 78147;
	#10 counter$count = 78148;
	#10 counter$count = 78149;
	#10 counter$count = 78150;
	#10 counter$count = 78151;
	#10 counter$count = 78152;
	#10 counter$count = 78153;
	#10 counter$count = 78154;
	#10 counter$count = 78155;
	#10 counter$count = 78156;
	#10 counter$count = 78157;
	#10 counter$count = 78158;
	#10 counter$count = 78159;
	#10 counter$count = 78160;
	#10 counter$count = 78161;
	#10 counter$count = 78162;
	#10 counter$count = 78163;
	#10 counter$count = 78164;
	#10 counter$count = 78165;
	#10 counter$count = 78166;
	#10 counter$count = 78167;
	#10 counter$count = 78168;
	#10 counter$count = 78169;
	#10 counter$count = 78170;
	#10 counter$count = 78171;
	#10 counter$count = 78172;
	#10 counter$count = 78173;
	#10 counter$count = 78174;
	#10 counter$count = 78175;
	#10 counter$count = 78176;
	#10 counter$count = 78177;
	#10 counter$count = 78178;
	#10 counter$count = 78179;
	#10 counter$count = 78180;
	#10 counter$count = 78181;
	#10 counter$count = 78182;
	#10 counter$count = 78183;
	#10 counter$count = 78184;
	#10 counter$count = 78185;
	#10 counter$count = 78186;
	#10 counter$count = 78187;
	#10 counter$count = 78188;
	#10 counter$count = 78189;
	#10 counter$count = 78190;
	#10 counter$count = 78191;
	#10 counter$count = 78192;
	#10 counter$count = 78193;
	#10 counter$count = 78194;
	#10 counter$count = 78195;
	#10 counter$count = 78196;
	#10 counter$count = 78197;
	#10 counter$count = 78198;
	#10 counter$count = 78199;
	#10 counter$count = 78200;
	#10 counter$count = 78201;
	#10 counter$count = 78202;
	#10 counter$count = 78203;
	#10 counter$count = 78204;
	#10 counter$count = 78205;
	#10 counter$count = 78206;
	#10 counter$count = 78207;
	#10 counter$count = 78208;
	#10 counter$count = 78209;
	#10 counter$count = 78210;
	#10 counter$count = 78211;
	#10 counter$count = 78212;
	#10 counter$count = 78213;
	#10 counter$count = 78214;
	#10 counter$count = 78215;
	#10 counter$count = 78216;
	#10 counter$count = 78217;
	#10 counter$count = 78218;
	#10 counter$count = 78219;
	#10 counter$count = 78220;
	#10 counter$count = 78221;
	#10 counter$count = 78222;
	#10 counter$count = 78223;
	#10 counter$count = 78224;
	#10 counter$count = 78225;
	#10 counter$count = 78226;
	#10 counter$count = 78227;
	#10 counter$count = 78228;
	#10 counter$count = 78229;
	#10 counter$count = 78230;
	#10 counter$count = 78231;
	#10 counter$count = 78232;
	#10 counter$count = 78233;
	#10 counter$count = 78234;
	#10 counter$count = 78235;
	#10 counter$count = 78236;
	#10 counter$count = 78237;
	#10 counter$count = 78238;
	#10 counter$count = 78239;
	#10 counter$count = 78240;
	#10 counter$count = 78241;
	#10 counter$count = 78242;
	#10 counter$count = 78243;
	#10 counter$count = 78244;
	#10 counter$count = 78245;
	#10 counter$count = 78246;
	#10 counter$count = 78247;
	#10 counter$count = 78248;
	#10 counter$count = 78249;
	#10 counter$count = 78250;
	#10 counter$count = 78251;
	#10 counter$count = 78252;
	#10 counter$count = 78253;
	#10 counter$count = 78254;
	#10 counter$count = 78255;
	#10 counter$count = 78256;
	#10 counter$count = 78257;
	#10 counter$count = 78258;
	#10 counter$count = 78259;
	#10 counter$count = 78260;
	#10 counter$count = 78261;
	#10 counter$count = 78262;
	#10 counter$count = 78263;
	#10 counter$count = 78264;
	#10 counter$count = 78265;
	#10 counter$count = 78266;
	#10 counter$count = 78267;
	#10 counter$count = 78268;
	#10 counter$count = 78269;
	#10 counter$count = 78270;
	#10 counter$count = 78271;
	#10 counter$count = 78272;
	#10 counter$count = 78273;
	#10 counter$count = 78274;
	#10 counter$count = 78275;
	#10 counter$count = 78276;
	#10 counter$count = 78277;
	#10 counter$count = 78278;
	#10 counter$count = 78279;
	#10 counter$count = 78280;
	#10 counter$count = 78281;
	#10 counter$count = 78282;
	#10 counter$count = 78283;
	#10 counter$count = 78284;
	#10 counter$count = 78285;
	#10 counter$count = 78286;
	#10 counter$count = 78287;
	#10 counter$count = 78288;
	#10 counter$count = 78289;
	#10 counter$count = 78290;
	#10 counter$count = 78291;
	#10 counter$count = 78292;
	#10 counter$count = 78293;
	#10 counter$count = 78294;
	#10 counter$count = 78295;
	#10 counter$count = 78296;
	#10 counter$count = 78297;
	#10 counter$count = 78298;
	#10 counter$count = 78299;
	#10 counter$count = 78300;
	#10 counter$count = 78301;
	#10 counter$count = 78302;
	#10 counter$count = 78303;
	#10 counter$count = 78304;
	#10 counter$count = 78305;
	#10 counter$count = 78306;
	#10 counter$count = 78307;
	#10 counter$count = 78308;
	#10 counter$count = 78309;
	#10 counter$count = 78310;
	#10 counter$count = 78311;
	#10 counter$count = 78312;
	#10 counter$count = 78313;
	#10 counter$count = 78314;
	#10 counter$count = 78315;
	#10 counter$count = 78316;
	#10 counter$count = 78317;
	#10 counter$count = 78318;
	#10 counter$count = 78319;
	#10 counter$count = 78320;
	#10 counter$count = 78321;
	#10 counter$count = 78322;
	#10 counter$count = 78323;
	#10 counter$count = 78324;
	#10 counter$count = 78325;
	#10 counter$count = 78326;
	#10 counter$count = 78327;
	#10 counter$count = 78328;
	#10 counter$count = 78329;
	#10 counter$count = 78330;
	#10 counter$count = 78331;
	#10 counter$count = 78332;
	#10 counter$count = 78333;
	#10 counter$count = 78334;
	#10 counter$count = 78335;
	#10 counter$count = 78336;
	#10 counter$count = 78337;
	#10 counter$count = 78338;
	#10 counter$count = 78339;
	#10 counter$count = 78340;
	#10 counter$count = 78341;
	#10 counter$count = 78342;
	#10 counter$count = 78343;
	#10 counter$count = 78344;
	#10 counter$count = 78345;
	#10 counter$count = 78346;
	#10 counter$count = 78347;
	#10 counter$count = 78348;
	#10 counter$count = 78349;
	#10 counter$count = 78350;
	#10 counter$count = 78351;
	#10 counter$count = 78352;
	#10 counter$count = 78353;
	#10 counter$count = 78354;
	#10 counter$count = 78355;
	#10 counter$count = 78356;
	#10 counter$count = 78357;
	#10 counter$count = 78358;
	#10 counter$count = 78359;
	#10 counter$count = 78360;
	#10 counter$count = 78361;
	#10 counter$count = 78362;
	#10 counter$count = 78363;
	#10 counter$count = 78364;
	#10 counter$count = 78365;
	#10 counter$count = 78366;
	#10 counter$count = 78367;
	#10 counter$count = 78368;
	#10 counter$count = 78369;
	#10 counter$count = 78370;
	#10 counter$count = 78371;
	#10 counter$count = 78372;
	#10 counter$count = 78373;
	#10 counter$count = 78374;
	#10 counter$count = 78375;
	#10 counter$count = 78376;
	#10 counter$count = 78377;
	#10 counter$count = 78378;
	#10 counter$count = 78379;
	#10 counter$count = 78380;
	#10 counter$count = 78381;
	#10 counter$count = 78382;
	#10 counter$count = 78383;
	#10 counter$count = 78384;
	#10 counter$count = 78385;
	#10 counter$count = 78386;
	#10 counter$count = 78387;
	#10 counter$count = 78388;
	#10 counter$count = 78389;
	#10 counter$count = 78390;
	#10 counter$count = 78391;
	#10 counter$count = 78392;
	#10 counter$count = 78393;
	#10 counter$count = 78394;
	#10 counter$count = 78395;
	#10 counter$count = 78396;
	#10 counter$count = 78397;
	#10 counter$count = 78398;
	#10 counter$count = 78399;
	#10 counter$count = 78400;
	#10 counter$count = 78401;
	#10 counter$count = 78402;
	#10 counter$count = 78403;
	#10 counter$count = 78404;
	#10 counter$count = 78405;
	#10 counter$count = 78406;
	#10 counter$count = 78407;
	#10 counter$count = 78408;
	#10 counter$count = 78409;
	#10 counter$count = 78410;
	#10 counter$count = 78411;
	#10 counter$count = 78412;
	#10 counter$count = 78413;
	#10 counter$count = 78414;
	#10 counter$count = 78415;
	#10 counter$count = 78416;
	#10 counter$count = 78417;
	#10 counter$count = 78418;
	#10 counter$count = 78419;
	#10 counter$count = 78420;
	#10 counter$count = 78421;
	#10 counter$count = 78422;
	#10 counter$count = 78423;
	#10 counter$count = 78424;
	#10 counter$count = 78425;
	#10 counter$count = 78426;
	#10 counter$count = 78427;
	#10 counter$count = 78428;
	#10 counter$count = 78429;
	#10 counter$count = 78430;
	#10 counter$count = 78431;
	#10 counter$count = 78432;
	#10 counter$count = 78433;
	#10 counter$count = 78434;
	#10 counter$count = 78435;
	#10 counter$count = 78436;
	#10 counter$count = 78437;
	#10 counter$count = 78438;
	#10 counter$count = 78439;
	#10 counter$count = 78440;
	#10 counter$count = 78441;
	#10 counter$count = 78442;
	#10 counter$count = 78443;
	#10 counter$count = 78444;
	#10 counter$count = 78445;
	#10 counter$count = 78446;
	#10 counter$count = 78447;
	#10 counter$count = 78448;
	#10 counter$count = 78449;
	#10 counter$count = 78450;
	#10 counter$count = 78451;
	#10 counter$count = 78452;
	#10 counter$count = 78453;
	#10 counter$count = 78454;
	#10 counter$count = 78455;
	#10 counter$count = 78456;
	#10 counter$count = 78457;
	#10 counter$count = 78458;
	#10 counter$count = 78459;
	#10 counter$count = 78460;
	#10 counter$count = 78461;
	#10 counter$count = 78462;
	#10 counter$count = 78463;
	#10 counter$count = 78464;
	#10 counter$count = 78465;
	#10 counter$count = 78466;
	#10 counter$count = 78467;
	#10 counter$count = 78468;
	#10 counter$count = 78469;
	#10 counter$count = 78470;
	#10 counter$count = 78471;
	#10 counter$count = 78472;
	#10 counter$count = 78473;
	#10 counter$count = 78474;
	#10 counter$count = 78475;
	#10 counter$count = 78476;
	#10 counter$count = 78477;
	#10 counter$count = 78478;
	#10 counter$count = 78479;
	#10 counter$count = 78480;
	#10 counter$count = 78481;
	#10 counter$count = 78482;
	#10 counter$count = 78483;
	#10 counter$count = 78484;
	#10 counter$count = 78485;
	#10 counter$count = 78486;
	#10 counter$count = 78487;
	#10 counter$count = 78488;
	#10 counter$count = 78489;
	#10 counter$count = 78490;
	#10 counter$count = 78491;
	#10 counter$count = 78492;
	#10 counter$count = 78493;
	#10 counter$count = 78494;
	#10 counter$count = 78495;
	#10 counter$count = 78496;
	#10 counter$count = 78497;
	#10 counter$count = 78498;
	#10 counter$count = 78499;
	#10 counter$count = 78500;
	#10 counter$count = 78501;
	#10 counter$count = 78502;
	#10 counter$count = 78503;
	#10 counter$count = 78504;
	#10 counter$count = 78505;
	#10 counter$count = 78506;
	#10 counter$count = 78507;
	#10 counter$count = 78508;
	#10 counter$count = 78509;
	#10 counter$count = 78510;
	#10 counter$count = 78511;
	#10 counter$count = 78512;
	#10 counter$count = 78513;
	#10 counter$count = 78514;
	#10 counter$count = 78515;
	#10 counter$count = 78516;
	#10 counter$count = 78517;
	#10 counter$count = 78518;
	#10 counter$count = 78519;
	#10 counter$count = 78520;
	#10 counter$count = 78521;
	#10 counter$count = 78522;
	#10 counter$count = 78523;
	#10 counter$count = 78524;
	#10 counter$count = 78525;
	#10 counter$count = 78526;
	#10 counter$count = 78527;
	#10 counter$count = 78528;
	#10 counter$count = 78529;
	#10 counter$count = 78530;
	#10 counter$count = 78531;
	#10 counter$count = 78532;
	#10 counter$count = 78533;
	#10 counter$count = 78534;
	#10 counter$count = 78535;
	#10 counter$count = 78536;
	#10 counter$count = 78537;
	#10 counter$count = 78538;
	#10 counter$count = 78539;
	#10 counter$count = 78540;
	#10 counter$count = 78541;
	#10 counter$count = 78542;
	#10 counter$count = 78543;
	#10 counter$count = 78544;
	#10 counter$count = 78545;
	#10 counter$count = 78546;
	#10 counter$count = 78547;
	#10 counter$count = 78548;
	#10 counter$count = 78549;
	#10 counter$count = 78550;
	#10 counter$count = 78551;
	#10 counter$count = 78552;
	#10 counter$count = 78553;
	#10 counter$count = 78554;
	#10 counter$count = 78555;
	#10 counter$count = 78556;
	#10 counter$count = 78557;
	#10 counter$count = 78558;
	#10 counter$count = 78559;
	#10 counter$count = 78560;
	#10 counter$count = 78561;
	#10 counter$count = 78562;
	#10 counter$count = 78563;
	#10 counter$count = 78564;
	#10 counter$count = 78565;
	#10 counter$count = 78566;
	#10 counter$count = 78567;
	#10 counter$count = 78568;
	#10 counter$count = 78569;
	#10 counter$count = 78570;
	#10 counter$count = 78571;
	#10 counter$count = 78572;
	#10 counter$count = 78573;
	#10 counter$count = 78574;
	#10 counter$count = 78575;
	#10 counter$count = 78576;
	#10 counter$count = 78577;
	#10 counter$count = 78578;
	#10 counter$count = 78579;
	#10 counter$count = 78580;
	#10 counter$count = 78581;
	#10 counter$count = 78582;
	#10 counter$count = 78583;
	#10 counter$count = 78584;
	#10 counter$count = 78585;
	#10 counter$count = 78586;
	#10 counter$count = 78587;
	#10 counter$count = 78588;
	#10 counter$count = 78589;
	#10 counter$count = 78590;
	#10 counter$count = 78591;
	#10 counter$count = 78592;
	#10 counter$count = 78593;
	#10 counter$count = 78594;
	#10 counter$count = 78595;
	#10 counter$count = 78596;
	#10 counter$count = 78597;
	#10 counter$count = 78598;
	#10 counter$count = 78599;
	#10 counter$count = 78600;
	#10 counter$count = 78601;
	#10 counter$count = 78602;
	#10 counter$count = 78603;
	#10 counter$count = 78604;
	#10 counter$count = 78605;
	#10 counter$count = 78606;
	#10 counter$count = 78607;
	#10 counter$count = 78608;
	#10 counter$count = 78609;
	#10 counter$count = 78610;
	#10 counter$count = 78611;
	#10 counter$count = 78612;
	#10 counter$count = 78613;
	#10 counter$count = 78614;
	#10 counter$count = 78615;
	#10 counter$count = 78616;
	#10 counter$count = 78617;
	#10 counter$count = 78618;
	#10 counter$count = 78619;
	#10 counter$count = 78620;
	#10 counter$count = 78621;
	#10 counter$count = 78622;
	#10 counter$count = 78623;
	#10 counter$count = 78624;
	#10 counter$count = 78625;
	#10 counter$count = 78626;
	#10 counter$count = 78627;
	#10 counter$count = 78628;
	#10 counter$count = 78629;
	#10 counter$count = 78630;
	#10 counter$count = 78631;
	#10 counter$count = 78632;
	#10 counter$count = 78633;
	#10 counter$count = 78634;
	#10 counter$count = 78635;
	#10 counter$count = 78636;
	#10 counter$count = 78637;
	#10 counter$count = 78638;
	#10 counter$count = 78639;
	#10 counter$count = 78640;
	#10 counter$count = 78641;
	#10 counter$count = 78642;
	#10 counter$count = 78643;
	#10 counter$count = 78644;
	#10 counter$count = 78645;
	#10 counter$count = 78646;
	#10 counter$count = 78647;
	#10 counter$count = 78648;
	#10 counter$count = 78649;
	#10 counter$count = 78650;
	#10 counter$count = 78651;
	#10 counter$count = 78652;
	#10 counter$count = 78653;
	#10 counter$count = 78654;
	#10 counter$count = 78655;
	#10 counter$count = 78656;
	#10 counter$count = 78657;
	#10 counter$count = 78658;
	#10 counter$count = 78659;
	#10 counter$count = 78660;
	#10 counter$count = 78661;
	#10 counter$count = 78662;
	#10 counter$count = 78663;
	#10 counter$count = 78664;
	#10 counter$count = 78665;
	#10 counter$count = 78666;
	#10 counter$count = 78667;
	#10 counter$count = 78668;
	#10 counter$count = 78669;
	#10 counter$count = 78670;
	#10 counter$count = 78671;
	#10 counter$count = 78672;
	#10 counter$count = 78673;
	#10 counter$count = 78674;
	#10 counter$count = 78675;
	#10 counter$count = 78676;
	#10 counter$count = 78677;
	#10 counter$count = 78678;
	#10 counter$count = 78679;
	#10 counter$count = 78680;
	#10 counter$count = 78681;
	#10 counter$count = 78682;
	#10 counter$count = 78683;
	#10 counter$count = 78684;
	#10 counter$count = 78685;
	#10 counter$count = 78686;
	#10 counter$count = 78687;
	#10 counter$count = 78688;
	#10 counter$count = 78689;
	#10 counter$count = 78690;
	#10 counter$count = 78691;
	#10 counter$count = 78692;
	#10 counter$count = 78693;
	#10 counter$count = 78694;
	#10 counter$count = 78695;
	#10 counter$count = 78696;
	#10 counter$count = 78697;
	#10 counter$count = 78698;
	#10 counter$count = 78699;
	#10 counter$count = 78700;
	#10 counter$count = 78701;
	#10 counter$count = 78702;
	#10 counter$count = 78703;
	#10 counter$count = 78704;
	#10 counter$count = 78705;
	#10 counter$count = 78706;
	#10 counter$count = 78707;
	#10 counter$count = 78708;
	#10 counter$count = 78709;
	#10 counter$count = 78710;
	#10 counter$count = 78711;
	#10 counter$count = 78712;
	#10 counter$count = 78713;
	#10 counter$count = 78714;
	#10 counter$count = 78715;
	#10 counter$count = 78716;
	#10 counter$count = 78717;
	#10 counter$count = 78718;
	#10 counter$count = 78719;
	#10 counter$count = 78720;
	#10 counter$count = 78721;
	#10 counter$count = 78722;
	#10 counter$count = 78723;
	#10 counter$count = 78724;
	#10 counter$count = 78725;
	#10 counter$count = 78726;
	#10 counter$count = 78727;
	#10 counter$count = 78728;
	#10 counter$count = 78729;
	#10 counter$count = 78730;
	#10 counter$count = 78731;
	#10 counter$count = 78732;
	#10 counter$count = 78733;
	#10 counter$count = 78734;
	#10 counter$count = 78735;
	#10 counter$count = 78736;
	#10 counter$count = 78737;
	#10 counter$count = 78738;
	#10 counter$count = 78739;
	#10 counter$count = 78740;
	#10 counter$count = 78741;
	#10 counter$count = 78742;
	#10 counter$count = 78743;
	#10 counter$count = 78744;
	#10 counter$count = 78745;
	#10 counter$count = 78746;
	#10 counter$count = 78747;
	#10 counter$count = 78748;
	#10 counter$count = 78749;
	#10 counter$count = 78750;
	#10 counter$count = 78751;
	#10 counter$count = 78752;
	#10 counter$count = 78753;
	#10 counter$count = 78754;
	#10 counter$count = 78755;
	#10 counter$count = 78756;
	#10 counter$count = 78757;
	#10 counter$count = 78758;
	#10 counter$count = 78759;
	#10 counter$count = 78760;
	#10 counter$count = 78761;
	#10 counter$count = 78762;
	#10 counter$count = 78763;
	#10 counter$count = 78764;
	#10 counter$count = 78765;
	#10 counter$count = 78766;
	#10 counter$count = 78767;
	#10 counter$count = 78768;
	#10 counter$count = 78769;
	#10 counter$count = 78770;
	#10 counter$count = 78771;
	#10 counter$count = 78772;
	#10 counter$count = 78773;
	#10 counter$count = 78774;
	#10 counter$count = 78775;
	#10 counter$count = 78776;
	#10 counter$count = 78777;
	#10 counter$count = 78778;
	#10 counter$count = 78779;
	#10 counter$count = 78780;
	#10 counter$count = 78781;
	#10 counter$count = 78782;
	#10 counter$count = 78783;
	#10 counter$count = 78784;
	#10 counter$count = 78785;
	#10 counter$count = 78786;
	#10 counter$count = 78787;
	#10 counter$count = 78788;
	#10 counter$count = 78789;
	#10 counter$count = 78790;
	#10 counter$count = 78791;
	#10 counter$count = 78792;
	#10 counter$count = 78793;
	#10 counter$count = 78794;
	#10 counter$count = 78795;
	#10 counter$count = 78796;
	#10 counter$count = 78797;
	#10 counter$count = 78798;
	#10 counter$count = 78799;
	#10 counter$count = 78800;
	#10 counter$count = 78801;
	#10 counter$count = 78802;
	#10 counter$count = 78803;
	#10 counter$count = 78804;
	#10 counter$count = 78805;
	#10 counter$count = 78806;
	#10 counter$count = 78807;
	#10 counter$count = 78808;
	#10 counter$count = 78809;
	#10 counter$count = 78810;
	#10 counter$count = 78811;
	#10 counter$count = 78812;
	#10 counter$count = 78813;
	#10 counter$count = 78814;
	#10 counter$count = 78815;
	#10 counter$count = 78816;
	#10 counter$count = 78817;
	#10 counter$count = 78818;
	#10 counter$count = 78819;
	#10 counter$count = 78820;
	#10 counter$count = 78821;
	#10 counter$count = 78822;
	#10 counter$count = 78823;
	#10 counter$count = 78824;
	#10 counter$count = 78825;
	#10 counter$count = 78826;
	#10 counter$count = 78827;
	#10 counter$count = 78828;
	#10 counter$count = 78829;
	#10 counter$count = 78830;
	#10 counter$count = 78831;
	#10 counter$count = 78832;
	#10 counter$count = 78833;
	#10 counter$count = 78834;
	#10 counter$count = 78835;
	#10 counter$count = 78836;
	#10 counter$count = 78837;
	#10 counter$count = 78838;
	#10 counter$count = 78839;
	#10 counter$count = 78840;
	#10 counter$count = 78841;
	#10 counter$count = 78842;
	#10 counter$count = 78843;
	#10 counter$count = 78844;
	#10 counter$count = 78845;
	#10 counter$count = 78846;
	#10 counter$count = 78847;
	#10 counter$count = 78848;
	#10 counter$count = 78849;
	#10 counter$count = 78850;
	#10 counter$count = 78851;
	#10 counter$count = 78852;
	#10 counter$count = 78853;
	#10 counter$count = 78854;
	#10 counter$count = 78855;
	#10 counter$count = 78856;
	#10 counter$count = 78857;
	#10 counter$count = 78858;
	#10 counter$count = 78859;
	#10 counter$count = 78860;
	#10 counter$count = 78861;
	#10 counter$count = 78862;
	#10 counter$count = 78863;
	#10 counter$count = 78864;
	#10 counter$count = 78865;
	#10 counter$count = 78866;
	#10 counter$count = 78867;
	#10 counter$count = 78868;
	#10 counter$count = 78869;
	#10 counter$count = 78870;
	#10 counter$count = 78871;
	#10 counter$count = 78872;
	#10 counter$count = 78873;
	#10 counter$count = 78874;
	#10 counter$count = 78875;
	#10 counter$count = 78876;
	#10 counter$count = 78877;
	#10 counter$count = 78878;
	#10 counter$count = 78879;
	#10 counter$count = 78880;
	#10 counter$count = 78881;
	#10 counter$count = 78882;
	#10 counter$count = 78883;
	#10 counter$count = 78884;
	#10 counter$count = 78885;
	#10 counter$count = 78886;
	#10 counter$count = 78887;
	#10 counter$count = 78888;
	#10 counter$count = 78889;
	#10 counter$count = 78890;
	#10 counter$count = 78891;
	#10 counter$count = 78892;
	#10 counter$count = 78893;
	#10 counter$count = 78894;
	#10 counter$count = 78895;
	#10 counter$count = 78896;
	#10 counter$count = 78897;
	#10 counter$count = 78898;
	#10 counter$count = 78899;
	#10 counter$count = 78900;
	#10 counter$count = 78901;
	#10 counter$count = 78902;
	#10 counter$count = 78903;
	#10 counter$count = 78904;
	#10 counter$count = 78905;
	#10 counter$count = 78906;
	#10 counter$count = 78907;
	#10 counter$count = 78908;
	#10 counter$count = 78909;
	#10 counter$count = 78910;
	#10 counter$count = 78911;
	#10 counter$count = 78912;
	#10 counter$count = 78913;
	#10 counter$count = 78914;
	#10 counter$count = 78915;
	#10 counter$count = 78916;
	#10 counter$count = 78917;
	#10 counter$count = 78918;
	#10 counter$count = 78919;
	#10 counter$count = 78920;
	#10 counter$count = 78921;
	#10 counter$count = 78922;
	#10 counter$count = 78923;
	#10 counter$count = 78924;
	#10 counter$count = 78925;
	#10 counter$count = 78926;
	#10 counter$count = 78927;
	#10 counter$count = 78928;
	#10 counter$count = 78929;
	#10 counter$count = 78930;
	#10 counter$count = 78931;
	#10 counter$count = 78932;
	#10 counter$count = 78933;
	#10 counter$count = 78934;
	#10 counter$count = 78935;
	#10 counter$count = 78936;
	#10 counter$count = 78937;
	#10 counter$count = 78938;
	#10 counter$count = 78939;
	#10 counter$count = 78940;
	#10 counter$count = 78941;
	#10 counter$count = 78942;
	#10 counter$count = 78943;
	#10 counter$count = 78944;
	#10 counter$count = 78945;
	#10 counter$count = 78946;
	#10 counter$count = 78947;
	#10 counter$count = 78948;
	#10 counter$count = 78949;
	#10 counter$count = 78950;
	#10 counter$count = 78951;
	#10 counter$count = 78952;
	#10 counter$count = 78953;
	#10 counter$count = 78954;
	#10 counter$count = 78955;
	#10 counter$count = 78956;
	#10 counter$count = 78957;
	#10 counter$count = 78958;
	#10 counter$count = 78959;
	#10 counter$count = 78960;
	#10 counter$count = 78961;
	#10 counter$count = 78962;
	#10 counter$count = 78963;
	#10 counter$count = 78964;
	#10 counter$count = 78965;
	#10 counter$count = 78966;
	#10 counter$count = 78967;
	#10 counter$count = 78968;
	#10 counter$count = 78969;
	#10 counter$count = 78970;
	#10 counter$count = 78971;
	#10 counter$count = 78972;
	#10 counter$count = 78973;
	#10 counter$count = 78974;
	#10 counter$count = 78975;
	#10 counter$count = 78976;
	#10 counter$count = 78977;
	#10 counter$count = 78978;
	#10 counter$count = 78979;
	#10 counter$count = 78980;
	#10 counter$count = 78981;
	#10 counter$count = 78982;
	#10 counter$count = 78983;
	#10 counter$count = 78984;
	#10 counter$count = 78985;
	#10 counter$count = 78986;
	#10 counter$count = 78987;
	#10 counter$count = 78988;
	#10 counter$count = 78989;
	#10 counter$count = 78990;
	#10 counter$count = 78991;
	#10 counter$count = 78992;
	#10 counter$count = 78993;
	#10 counter$count = 78994;
	#10 counter$count = 78995;
	#10 counter$count = 78996;
	#10 counter$count = 78997;
	#10 counter$count = 78998;
	#10 counter$count = 78999;
	#10 counter$count = 79000;
	#10 counter$count = 79001;
	#10 counter$count = 79002;
	#10 counter$count = 79003;
	#10 counter$count = 79004;
	#10 counter$count = 79005;
	#10 counter$count = 79006;
	#10 counter$count = 79007;
	#10 counter$count = 79008;
	#10 counter$count = 79009;
	#10 counter$count = 79010;
	#10 counter$count = 79011;
	#10 counter$count = 79012;
	#10 counter$count = 79013;
	#10 counter$count = 79014;
	#10 counter$count = 79015;
	#10 counter$count = 79016;
	#10 counter$count = 79017;
	#10 counter$count = 79018;
	#10 counter$count = 79019;
	#10 counter$count = 79020;
	#10 counter$count = 79021;
	#10 counter$count = 79022;
	#10 counter$count = 79023;
	#10 counter$count = 79024;
	#10 counter$count = 79025;
	#10 counter$count = 79026;
	#10 counter$count = 79027;
	#10 counter$count = 79028;
	#10 counter$count = 79029;
	#10 counter$count = 79030;
	#10 counter$count = 79031;
	#10 counter$count = 79032;
	#10 counter$count = 79033;
	#10 counter$count = 79034;
	#10 counter$count = 79035;
	#10 counter$count = 79036;
	#10 counter$count = 79037;
	#10 counter$count = 79038;
	#10 counter$count = 79039;
	#10 counter$count = 79040;
	#10 counter$count = 79041;
	#10 counter$count = 79042;
	#10 counter$count = 79043;
	#10 counter$count = 79044;
	#10 counter$count = 79045;
	#10 counter$count = 79046;
	#10 counter$count = 79047;
	#10 counter$count = 79048;
	#10 counter$count = 79049;
	#10 counter$count = 79050;
	#10 counter$count = 79051;
	#10 counter$count = 79052;
	#10 counter$count = 79053;
	#10 counter$count = 79054;
	#10 counter$count = 79055;
	#10 counter$count = 79056;
	#10 counter$count = 79057;
	#10 counter$count = 79058;
	#10 counter$count = 79059;
	#10 counter$count = 79060;
	#10 counter$count = 79061;
	#10 counter$count = 79062;
	#10 counter$count = 79063;
	#10 counter$count = 79064;
	#10 counter$count = 79065;
	#10 counter$count = 79066;
	#10 counter$count = 79067;
	#10 counter$count = 79068;
	#10 counter$count = 79069;
	#10 counter$count = 79070;
	#10 counter$count = 79071;
	#10 counter$count = 79072;
	#10 counter$count = 79073;
	#10 counter$count = 79074;
	#10 counter$count = 79075;
	#10 counter$count = 79076;
	#10 counter$count = 79077;
	#10 counter$count = 79078;
	#10 counter$count = 79079;
	#10 counter$count = 79080;
	#10 counter$count = 79081;
	#10 counter$count = 79082;
	#10 counter$count = 79083;
	#10 counter$count = 79084;
	#10 counter$count = 79085;
	#10 counter$count = 79086;
	#10 counter$count = 79087;
	#10 counter$count = 79088;
	#10 counter$count = 79089;
	#10 counter$count = 79090;
	#10 counter$count = 79091;
	#10 counter$count = 79092;
	#10 counter$count = 79093;
	#10 counter$count = 79094;
	#10 counter$count = 79095;
	#10 counter$count = 79096;
	#10 counter$count = 79097;
	#10 counter$count = 79098;
	#10 counter$count = 79099;
	#10 counter$count = 79100;
	#10 counter$count = 79101;
	#10 counter$count = 79102;
	#10 counter$count = 79103;
	#10 counter$count = 79104;
	#10 counter$count = 79105;
	#10 counter$count = 79106;
	#10 counter$count = 79107;
	#10 counter$count = 79108;
	#10 counter$count = 79109;
	#10 counter$count = 79110;
	#10 counter$count = 79111;
	#10 counter$count = 79112;
	#10 counter$count = 79113;
	#10 counter$count = 79114;
	#10 counter$count = 79115;
	#10 counter$count = 79116;
	#10 counter$count = 79117;
	#10 counter$count = 79118;
	#10 counter$count = 79119;
	#10 counter$count = 79120;
	#10 counter$count = 79121;
	#10 counter$count = 79122;
	#10 counter$count = 79123;
	#10 counter$count = 79124;
	#10 counter$count = 79125;
	#10 counter$count = 79126;
	#10 counter$count = 79127;
	#10 counter$count = 79128;
	#10 counter$count = 79129;
	#10 counter$count = 79130;
	#10 counter$count = 79131;
	#10 counter$count = 79132;
	#10 counter$count = 79133;
	#10 counter$count = 79134;
	#10 counter$count = 79135;
	#10 counter$count = 79136;
	#10 counter$count = 79137;
	#10 counter$count = 79138;
	#10 counter$count = 79139;
	#10 counter$count = 79140;
	#10 counter$count = 79141;
	#10 counter$count = 79142;
	#10 counter$count = 79143;
	#10 counter$count = 79144;
	#10 counter$count = 79145;
	#10 counter$count = 79146;
	#10 counter$count = 79147;
	#10 counter$count = 79148;
	#10 counter$count = 79149;
	#10 counter$count = 79150;
	#10 counter$count = 79151;
	#10 counter$count = 79152;
	#10 counter$count = 79153;
	#10 counter$count = 79154;
	#10 counter$count = 79155;
	#10 counter$count = 79156;
	#10 counter$count = 79157;
	#10 counter$count = 79158;
	#10 counter$count = 79159;
	#10 counter$count = 79160;
	#10 counter$count = 79161;
	#10 counter$count = 79162;
	#10 counter$count = 79163;
	#10 counter$count = 79164;
	#10 counter$count = 79165;
	#10 counter$count = 79166;
	#10 counter$count = 79167;
	#10 counter$count = 79168;
	#10 counter$count = 79169;
	#10 counter$count = 79170;
	#10 counter$count = 79171;
	#10 counter$count = 79172;
	#10 counter$count = 79173;
	#10 counter$count = 79174;
	#10 counter$count = 79175;
	#10 counter$count = 79176;
	#10 counter$count = 79177;
	#10 counter$count = 79178;
	#10 counter$count = 79179;
	#10 counter$count = 79180;
	#10 counter$count = 79181;
	#10 counter$count = 79182;
	#10 counter$count = 79183;
	#10 counter$count = 79184;
	#10 counter$count = 79185;
	#10 counter$count = 79186;
	#10 counter$count = 79187;
	#10 counter$count = 79188;
	#10 counter$count = 79189;
	#10 counter$count = 79190;
	#10 counter$count = 79191;
	#10 counter$count = 79192;
	#10 counter$count = 79193;
	#10 counter$count = 79194;
	#10 counter$count = 79195;
	#10 counter$count = 79196;
	#10 counter$count = 79197;
	#10 counter$count = 79198;
	#10 counter$count = 79199;
	#10 counter$count = 79200;
	#10 counter$count = 79201;
	#10 counter$count = 79202;
	#10 counter$count = 79203;
	#10 counter$count = 79204;
	#10 counter$count = 79205;
	#10 counter$count = 79206;
	#10 counter$count = 79207;
	#10 counter$count = 79208;
	#10 counter$count = 79209;
	#10 counter$count = 79210;
	#10 counter$count = 79211;
	#10 counter$count = 79212;
	#10 counter$count = 79213;
	#10 counter$count = 79214;
	#10 counter$count = 79215;
	#10 counter$count = 79216;
	#10 counter$count = 79217;
	#10 counter$count = 79218;
	#10 counter$count = 79219;
	#10 counter$count = 79220;
	#10 counter$count = 79221;
	#10 counter$count = 79222;
	#10 counter$count = 79223;
	#10 counter$count = 79224;
	#10 counter$count = 79225;
	#10 counter$count = 79226;
	#10 counter$count = 79227;
	#10 counter$count = 79228;
	#10 counter$count = 79229;
	#10 counter$count = 79230;
	#10 counter$count = 79231;
	#10 counter$count = 79232;
	#10 counter$count = 79233;
	#10 counter$count = 79234;
	#10 counter$count = 79235;
	#10 counter$count = 79236;
	#10 counter$count = 79237;
	#10 counter$count = 79238;
	#10 counter$count = 79239;
	#10 counter$count = 79240;
	#10 counter$count = 79241;
	#10 counter$count = 79242;
	#10 counter$count = 79243;
	#10 counter$count = 79244;
	#10 counter$count = 79245;
	#10 counter$count = 79246;
	#10 counter$count = 79247;
	#10 counter$count = 79248;
	#10 counter$count = 79249;
	#10 counter$count = 79250;
	#10 counter$count = 79251;
	#10 counter$count = 79252;
	#10 counter$count = 79253;
	#10 counter$count = 79254;
	#10 counter$count = 79255;
	#10 counter$count = 79256;
	#10 counter$count = 79257;
	#10 counter$count = 79258;
	#10 counter$count = 79259;
	#10 counter$count = 79260;
	#10 counter$count = 79261;
	#10 counter$count = 79262;
	#10 counter$count = 79263;
	#10 counter$count = 79264;
	#10 counter$count = 79265;
	#10 counter$count = 79266;
	#10 counter$count = 79267;
	#10 counter$count = 79268;
	#10 counter$count = 79269;
	#10 counter$count = 79270;
	#10 counter$count = 79271;
	#10 counter$count = 79272;
	#10 counter$count = 79273;
	#10 counter$count = 79274;
	#10 counter$count = 79275;
	#10 counter$count = 79276;
	#10 counter$count = 79277;
	#10 counter$count = 79278;
	#10 counter$count = 79279;
	#10 counter$count = 79280;
	#10 counter$count = 79281;
	#10 counter$count = 79282;
	#10 counter$count = 79283;
	#10 counter$count = 79284;
	#10 counter$count = 79285;
	#10 counter$count = 79286;
	#10 counter$count = 79287;
	#10 counter$count = 79288;
	#10 counter$count = 79289;
	#10 counter$count = 79290;
	#10 counter$count = 79291;
	#10 counter$count = 79292;
	#10 counter$count = 79293;
	#10 counter$count = 79294;
	#10 counter$count = 79295;
	#10 counter$count = 79296;
	#10 counter$count = 79297;
	#10 counter$count = 79298;
	#10 counter$count = 79299;
	#10 counter$count = 79300;
	#10 counter$count = 79301;
	#10 counter$count = 79302;
	#10 counter$count = 79303;
	#10 counter$count = 79304;
	#10 counter$count = 79305;
	#10 counter$count = 79306;
	#10 counter$count = 79307;
	#10 counter$count = 79308;
	#10 counter$count = 79309;
	#10 counter$count = 79310;
	#10 counter$count = 79311;
	#10 counter$count = 79312;
	#10 counter$count = 79313;
	#10 counter$count = 79314;
	#10 counter$count = 79315;
	#10 counter$count = 79316;
	#10 counter$count = 79317;
	#10 counter$count = 79318;
	#10 counter$count = 79319;
	#10 counter$count = 79320;
	#10 counter$count = 79321;
	#10 counter$count = 79322;
	#10 counter$count = 79323;
	#10 counter$count = 79324;
	#10 counter$count = 79325;
	#10 counter$count = 79326;
	#10 counter$count = 79327;
	#10 counter$count = 79328;
	#10 counter$count = 79329;
	#10 counter$count = 79330;
	#10 counter$count = 79331;
	#10 counter$count = 79332;
	#10 counter$count = 79333;
	#10 counter$count = 79334;
	#10 counter$count = 79335;
	#10 counter$count = 79336;
	#10 counter$count = 79337;
	#10 counter$count = 79338;
	#10 counter$count = 79339;
	#10 counter$count = 79340;
	#10 counter$count = 79341;
	#10 counter$count = 79342;
	#10 counter$count = 79343;
	#10 counter$count = 79344;
	#10 counter$count = 79345;
	#10 counter$count = 79346;
	#10 counter$count = 79347;
	#10 counter$count = 79348;
	#10 counter$count = 79349;
	#10 counter$count = 79350;
	#10 counter$count = 79351;
	#10 counter$count = 79352;
	#10 counter$count = 79353;
	#10 counter$count = 79354;
	#10 counter$count = 79355;
	#10 counter$count = 79356;
	#10 counter$count = 79357;
	#10 counter$count = 79358;
	#10 counter$count = 79359;
	#10 counter$count = 79360;
	#10 counter$count = 79361;
	#10 counter$count = 79362;
	#10 counter$count = 79363;
	#10 counter$count = 79364;
	#10 counter$count = 79365;
	#10 counter$count = 79366;
	#10 counter$count = 79367;
	#10 counter$count = 79368;
	#10 counter$count = 79369;
	#10 counter$count = 79370;
	#10 counter$count = 79371;
	#10 counter$count = 79372;
	#10 counter$count = 79373;
	#10 counter$count = 79374;
	#10 counter$count = 79375;
	#10 counter$count = 79376;
	#10 counter$count = 79377;
	#10 counter$count = 79378;
	#10 counter$count = 79379;
	#10 counter$count = 79380;
	#10 counter$count = 79381;
	#10 counter$count = 79382;
	#10 counter$count = 79383;
	#10 counter$count = 79384;
	#10 counter$count = 79385;
	#10 counter$count = 79386;
	#10 counter$count = 79387;
	#10 counter$count = 79388;
	#10 counter$count = 79389;
	#10 counter$count = 79390;
	#10 counter$count = 79391;
	#10 counter$count = 79392;
	#10 counter$count = 79393;
	#10 counter$count = 79394;
	#10 counter$count = 79395;
	#10 counter$count = 79396;
	#10 counter$count = 79397;
	#10 counter$count = 79398;
	#10 counter$count = 79399;
	#10 counter$count = 79400;
	#10 counter$count = 79401;
	#10 counter$count = 79402;
	#10 counter$count = 79403;
	#10 counter$count = 79404;
	#10 counter$count = 79405;
	#10 counter$count = 79406;
	#10 counter$count = 79407;
	#10 counter$count = 79408;
	#10 counter$count = 79409;
	#10 counter$count = 79410;
	#10 counter$count = 79411;
	#10 counter$count = 79412;
	#10 counter$count = 79413;
	#10 counter$count = 79414;
	#10 counter$count = 79415;
	#10 counter$count = 79416;
	#10 counter$count = 79417;
	#10 counter$count = 79418;
	#10 counter$count = 79419;
	#10 counter$count = 79420;
	#10 counter$count = 79421;
	#10 counter$count = 79422;
	#10 counter$count = 79423;
	#10 counter$count = 79424;
	#10 counter$count = 79425;
	#10 counter$count = 79426;
	#10 counter$count = 79427;
	#10 counter$count = 79428;
	#10 counter$count = 79429;
	#10 counter$count = 79430;
	#10 counter$count = 79431;
	#10 counter$count = 79432;
	#10 counter$count = 79433;
	#10 counter$count = 79434;
	#10 counter$count = 79435;
	#10 counter$count = 79436;
	#10 counter$count = 79437;
	#10 counter$count = 79438;
	#10 counter$count = 79439;
	#10 counter$count = 79440;
	#10 counter$count = 79441;
	#10 counter$count = 79442;
	#10 counter$count = 79443;
	#10 counter$count = 79444;
	#10 counter$count = 79445;
	#10 counter$count = 79446;
	#10 counter$count = 79447;
	#10 counter$count = 79448;
	#10 counter$count = 79449;
	#10 counter$count = 79450;
	#10 counter$count = 79451;
	#10 counter$count = 79452;
	#10 counter$count = 79453;
	#10 counter$count = 79454;
	#10 counter$count = 79455;
	#10 counter$count = 79456;
	#10 counter$count = 79457;
	#10 counter$count = 79458;
	#10 counter$count = 79459;
	#10 counter$count = 79460;
	#10 counter$count = 79461;
	#10 counter$count = 79462;
	#10 counter$count = 79463;
	#10 counter$count = 79464;
	#10 counter$count = 79465;
	#10 counter$count = 79466;
	#10 counter$count = 79467;
	#10 counter$count = 79468;
	#10 counter$count = 79469;
	#10 counter$count = 79470;
	#10 counter$count = 79471;
	#10 counter$count = 79472;
	#10 counter$count = 79473;
	#10 counter$count = 79474;
	#10 counter$count = 79475;
	#10 counter$count = 79476;
	#10 counter$count = 79477;
	#10 counter$count = 79478;
	#10 counter$count = 79479;
	#10 counter$count = 79480;
	#10 counter$count = 79481;
	#10 counter$count = 79482;
	#10 counter$count = 79483;
	#10 counter$count = 79484;
	#10 counter$count = 79485;
	#10 counter$count = 79486;
	#10 counter$count = 79487;
	#10 counter$count = 79488;
	#10 counter$count = 79489;
	#10 counter$count = 79490;
	#10 counter$count = 79491;
	#10 counter$count = 79492;
	#10 counter$count = 79493;
	#10 counter$count = 79494;
	#10 counter$count = 79495;
	#10 counter$count = 79496;
	#10 counter$count = 79497;
	#10 counter$count = 79498;
	#10 counter$count = 79499;
	#10 counter$count = 79500;
	#10 counter$count = 79501;
	#10 counter$count = 79502;
	#10 counter$count = 79503;
	#10 counter$count = 79504;
	#10 counter$count = 79505;
	#10 counter$count = 79506;
	#10 counter$count = 79507;
	#10 counter$count = 79508;
	#10 counter$count = 79509;
	#10 counter$count = 79510;
	#10 counter$count = 79511;
	#10 counter$count = 79512;
	#10 counter$count = 79513;
	#10 counter$count = 79514;
	#10 counter$count = 79515;
	#10 counter$count = 79516;
	#10 counter$count = 79517;
	#10 counter$count = 79518;
	#10 counter$count = 79519;
	#10 counter$count = 79520;
	#10 counter$count = 79521;
	#10 counter$count = 79522;
	#10 counter$count = 79523;
	#10 counter$count = 79524;
	#10 counter$count = 79525;
	#10 counter$count = 79526;
	#10 counter$count = 79527;
	#10 counter$count = 79528;
	#10 counter$count = 79529;
	#10 counter$count = 79530;
	#10 counter$count = 79531;
	#10 counter$count = 79532;
	#10 counter$count = 79533;
	#10 counter$count = 79534;
	#10 counter$count = 79535;
	#10 counter$count = 79536;
	#10 counter$count = 79537;
	#10 counter$count = 79538;
	#10 counter$count = 79539;
	#10 counter$count = 79540;
	#10 counter$count = 79541;
	#10 counter$count = 79542;
	#10 counter$count = 79543;
	#10 counter$count = 79544;
	#10 counter$count = 79545;
	#10 counter$count = 79546;
	#10 counter$count = 79547;
	#10 counter$count = 79548;
	#10 counter$count = 79549;
	#10 counter$count = 79550;
	#10 counter$count = 79551;
	#10 counter$count = 79552;
	#10 counter$count = 79553;
	#10 counter$count = 79554;
	#10 counter$count = 79555;
	#10 counter$count = 79556;
	#10 counter$count = 79557;
	#10 counter$count = 79558;
	#10 counter$count = 79559;
	#10 counter$count = 79560;
	#10 counter$count = 79561;
	#10 counter$count = 79562;
	#10 counter$count = 79563;
	#10 counter$count = 79564;
	#10 counter$count = 79565;
	#10 counter$count = 79566;
	#10 counter$count = 79567;
	#10 counter$count = 79568;
	#10 counter$count = 79569;
	#10 counter$count = 79570;
	#10 counter$count = 79571;
	#10 counter$count = 79572;
	#10 counter$count = 79573;
	#10 counter$count = 79574;
	#10 counter$count = 79575;
	#10 counter$count = 79576;
	#10 counter$count = 79577;
	#10 counter$count = 79578;
	#10 counter$count = 79579;
	#10 counter$count = 79580;
	#10 counter$count = 79581;
	#10 counter$count = 79582;
	#10 counter$count = 79583;
	#10 counter$count = 79584;
	#10 counter$count = 79585;
	#10 counter$count = 79586;
	#10 counter$count = 79587;
	#10 counter$count = 79588;
	#10 counter$count = 79589;
	#10 counter$count = 79590;
	#10 counter$count = 79591;
	#10 counter$count = 79592;
	#10 counter$count = 79593;
	#10 counter$count = 79594;
	#10 counter$count = 79595;
	#10 counter$count = 79596;
	#10 counter$count = 79597;
	#10 counter$count = 79598;
	#10 counter$count = 79599;
	#10 counter$count = 79600;
	#10 counter$count = 79601;
	#10 counter$count = 79602;
	#10 counter$count = 79603;
	#10 counter$count = 79604;
	#10 counter$count = 79605;
	#10 counter$count = 79606;
	#10 counter$count = 79607;
	#10 counter$count = 79608;
	#10 counter$count = 79609;
	#10 counter$count = 79610;
	#10 counter$count = 79611;
	#10 counter$count = 79612;
	#10 counter$count = 79613;
	#10 counter$count = 79614;
	#10 counter$count = 79615;
	#10 counter$count = 79616;
	#10 counter$count = 79617;
	#10 counter$count = 79618;
	#10 counter$count = 79619;
	#10 counter$count = 79620;
	#10 counter$count = 79621;
	#10 counter$count = 79622;
	#10 counter$count = 79623;
	#10 counter$count = 79624;
	#10 counter$count = 79625;
	#10 counter$count = 79626;
	#10 counter$count = 79627;
	#10 counter$count = 79628;
	#10 counter$count = 79629;
	#10 counter$count = 79630;
	#10 counter$count = 79631;
	#10 counter$count = 79632;
	#10 counter$count = 79633;
	#10 counter$count = 79634;
	#10 counter$count = 79635;
	#10 counter$count = 79636;
	#10 counter$count = 79637;
	#10 counter$count = 79638;
	#10 counter$count = 79639;
	#10 counter$count = 79640;
	#10 counter$count = 79641;
	#10 counter$count = 79642;
	#10 counter$count = 79643;
	#10 counter$count = 79644;
	#10 counter$count = 79645;
	#10 counter$count = 79646;
	#10 counter$count = 79647;
	#10 counter$count = 79648;
	#10 counter$count = 79649;
	#10 counter$count = 79650;
	#10 counter$count = 79651;
	#10 counter$count = 79652;
	#10 counter$count = 79653;
	#10 counter$count = 79654;
	#10 counter$count = 79655;
	#10 counter$count = 79656;
	#10 counter$count = 79657;
	#10 counter$count = 79658;
	#10 counter$count = 79659;
	#10 counter$count = 79660;
	#10 counter$count = 79661;
	#10 counter$count = 79662;
	#10 counter$count = 79663;
	#10 counter$count = 79664;
	#10 counter$count = 79665;
	#10 counter$count = 79666;
	#10 counter$count = 79667;
	#10 counter$count = 79668;
	#10 counter$count = 79669;
	#10 counter$count = 79670;
	#10 counter$count = 79671;
	#10 counter$count = 79672;
	#10 counter$count = 79673;
	#10 counter$count = 79674;
	#10 counter$count = 79675;
	#10 counter$count = 79676;
	#10 counter$count = 79677;
	#10 counter$count = 79678;
	#10 counter$count = 79679;
	#10 counter$count = 79680;
	#10 counter$count = 79681;
	#10 counter$count = 79682;
	#10 counter$count = 79683;
	#10 counter$count = 79684;
	#10 counter$count = 79685;
	#10 counter$count = 79686;
	#10 counter$count = 79687;
	#10 counter$count = 79688;
	#10 counter$count = 79689;
	#10 counter$count = 79690;
	#10 counter$count = 79691;
	#10 counter$count = 79692;
	#10 counter$count = 79693;
	#10 counter$count = 79694;
	#10 counter$count = 79695;
	#10 counter$count = 79696;
	#10 counter$count = 79697;
	#10 counter$count = 79698;
	#10 counter$count = 79699;
	#10 counter$count = 79700;
	#10 counter$count = 79701;
	#10 counter$count = 79702;
	#10 counter$count = 79703;
	#10 counter$count = 79704;
	#10 counter$count = 79705;
	#10 counter$count = 79706;
	#10 counter$count = 79707;
	#10 counter$count = 79708;
	#10 counter$count = 79709;
	#10 counter$count = 79710;
	#10 counter$count = 79711;
	#10 counter$count = 79712;
	#10 counter$count = 79713;
	#10 counter$count = 79714;
	#10 counter$count = 79715;
	#10 counter$count = 79716;
	#10 counter$count = 79717;
	#10 counter$count = 79718;
	#10 counter$count = 79719;
	#10 counter$count = 79720;
	#10 counter$count = 79721;
	#10 counter$count = 79722;
	#10 counter$count = 79723;
	#10 counter$count = 79724;
	#10 counter$count = 79725;
	#10 counter$count = 79726;
	#10 counter$count = 79727;
	#10 counter$count = 79728;
	#10 counter$count = 79729;
	#10 counter$count = 79730;
	#10 counter$count = 79731;
	#10 counter$count = 79732;
	#10 counter$count = 79733;
	#10 counter$count = 79734;
	#10 counter$count = 79735;
	#10 counter$count = 79736;
	#10 counter$count = 79737;
	#10 counter$count = 79738;
	#10 counter$count = 79739;
	#10 counter$count = 79740;
	#10 counter$count = 79741;
	#10 counter$count = 79742;
	#10 counter$count = 79743;
	#10 counter$count = 79744;
	#10 counter$count = 79745;
	#10 counter$count = 79746;
	#10 counter$count = 79747;
	#10 counter$count = 79748;
	#10 counter$count = 79749;
	#10 counter$count = 79750;
	#10 counter$count = 79751;
	#10 counter$count = 79752;
	#10 counter$count = 79753;
	#10 counter$count = 79754;
	#10 counter$count = 79755;
	#10 counter$count = 79756;
	#10 counter$count = 79757;
	#10 counter$count = 79758;
	#10 counter$count = 79759;
	#10 counter$count = 79760;
	#10 counter$count = 79761;
	#10 counter$count = 79762;
	#10 counter$count = 79763;
	#10 counter$count = 79764;
	#10 counter$count = 79765;
	#10 counter$count = 79766;
	#10 counter$count = 79767;
	#10 counter$count = 79768;
	#10 counter$count = 79769;
	#10 counter$count = 79770;
	#10 counter$count = 79771;
	#10 counter$count = 79772;
	#10 counter$count = 79773;
	#10 counter$count = 79774;
	#10 counter$count = 79775;
	#10 counter$count = 79776;
	#10 counter$count = 79777;
	#10 counter$count = 79778;
	#10 counter$count = 79779;
	#10 counter$count = 79780;
	#10 counter$count = 79781;
	#10 counter$count = 79782;
	#10 counter$count = 79783;
	#10 counter$count = 79784;
	#10 counter$count = 79785;
	#10 counter$count = 79786;
	#10 counter$count = 79787;
	#10 counter$count = 79788;
	#10 counter$count = 79789;
	#10 counter$count = 79790;
	#10 counter$count = 79791;
	#10 counter$count = 79792;
	#10 counter$count = 79793;
	#10 counter$count = 79794;
	#10 counter$count = 79795;
	#10 counter$count = 79796;
	#10 counter$count = 79797;
	#10 counter$count = 79798;
	#10 counter$count = 79799;
	#10 counter$count = 79800;
	#10 counter$count = 79801;
	#10 counter$count = 79802;
	#10 counter$count = 79803;
	#10 counter$count = 79804;
	#10 counter$count = 79805;
	#10 counter$count = 79806;
	#10 counter$count = 79807;
	#10 counter$count = 79808;
	#10 counter$count = 79809;
	#10 counter$count = 79810;
	#10 counter$count = 79811;
	#10 counter$count = 79812;
	#10 counter$count = 79813;
	#10 counter$count = 79814;
	#10 counter$count = 79815;
	#10 counter$count = 79816;
	#10 counter$count = 79817;
	#10 counter$count = 79818;
	#10 counter$count = 79819;
	#10 counter$count = 79820;
	#10 counter$count = 79821;
	#10 counter$count = 79822;
	#10 counter$count = 79823;
	#10 counter$count = 79824;
	#10 counter$count = 79825;
	#10 counter$count = 79826;
	#10 counter$count = 79827;
	#10 counter$count = 79828;
	#10 counter$count = 79829;
	#10 counter$count = 79830;
	#10 counter$count = 79831;
	#10 counter$count = 79832;
	#10 counter$count = 79833;
	#10 counter$count = 79834;
	#10 counter$count = 79835;
	#10 counter$count = 79836;
	#10 counter$count = 79837;
	#10 counter$count = 79838;
	#10 counter$count = 79839;
	#10 counter$count = 79840;
	#10 counter$count = 79841;
	#10 counter$count = 79842;
	#10 counter$count = 79843;
	#10 counter$count = 79844;
	#10 counter$count = 79845;
	#10 counter$count = 79846;
	#10 counter$count = 79847;
	#10 counter$count = 79848;
	#10 counter$count = 79849;
	#10 counter$count = 79850;
	#10 counter$count = 79851;
	#10 counter$count = 79852;
	#10 counter$count = 79853;
	#10 counter$count = 79854;
	#10 counter$count = 79855;
	#10 counter$count = 79856;
	#10 counter$count = 79857;
	#10 counter$count = 79858;
	#10 counter$count = 79859;
	#10 counter$count = 79860;
	#10 counter$count = 79861;
	#10 counter$count = 79862;
	#10 counter$count = 79863;
	#10 counter$count = 79864;
	#10 counter$count = 79865;
	#10 counter$count = 79866;
	#10 counter$count = 79867;
	#10 counter$count = 79868;
	#10 counter$count = 79869;
	#10 counter$count = 79870;
	#10 counter$count = 79871;
	#10 counter$count = 79872;
	#10 counter$count = 79873;
	#10 counter$count = 79874;
	#10 counter$count = 79875;
	#10 counter$count = 79876;
	#10 counter$count = 79877;
	#10 counter$count = 79878;
	#10 counter$count = 79879;
	#10 counter$count = 79880;
	#10 counter$count = 79881;
	#10 counter$count = 79882;
	#10 counter$count = 79883;
	#10 counter$count = 79884;
	#10 counter$count = 79885;
	#10 counter$count = 79886;
	#10 counter$count = 79887;
	#10 counter$count = 79888;
	#10 counter$count = 79889;
	#10 counter$count = 79890;
	#10 counter$count = 79891;
	#10 counter$count = 79892;
	#10 counter$count = 79893;
	#10 counter$count = 79894;
	#10 counter$count = 79895;
	#10 counter$count = 79896;
	#10 counter$count = 79897;
	#10 counter$count = 79898;
	#10 counter$count = 79899;
	#10 counter$count = 79900;
	#10 counter$count = 79901;
	#10 counter$count = 79902;
	#10 counter$count = 79903;
	#10 counter$count = 79904;
	#10 counter$count = 79905;
	#10 counter$count = 79906;
	#10 counter$count = 79907;
	#10 counter$count = 79908;
	#10 counter$count = 79909;
	#10 counter$count = 79910;
	#10 counter$count = 79911;
	#10 counter$count = 79912;
	#10 counter$count = 79913;
	#10 counter$count = 79914;
	#10 counter$count = 79915;
	#10 counter$count = 79916;
	#10 counter$count = 79917;
	#10 counter$count = 79918;
	#10 counter$count = 79919;
	#10 counter$count = 79920;
	#10 counter$count = 79921;
	#10 counter$count = 79922;
	#10 counter$count = 79923;
	#10 counter$count = 79924;
	#10 counter$count = 79925;
	#10 counter$count = 79926;
	#10 counter$count = 79927;
	#10 counter$count = 79928;
	#10 counter$count = 79929;
	#10 counter$count = 79930;
	#10 counter$count = 79931;
	#10 counter$count = 79932;
	#10 counter$count = 79933;
	#10 counter$count = 79934;
	#10 counter$count = 79935;
	#10 counter$count = 79936;
	#10 counter$count = 79937;
	#10 counter$count = 79938;
	#10 counter$count = 79939;
	#10 counter$count = 79940;
	#10 counter$count = 79941;
	#10 counter$count = 79942;
	#10 counter$count = 79943;
	#10 counter$count = 79944;
	#10 counter$count = 79945;
	#10 counter$count = 79946;
	#10 counter$count = 79947;
	#10 counter$count = 79948;
	#10 counter$count = 79949;
	#10 counter$count = 79950;
	#10 counter$count = 79951;
	#10 counter$count = 79952;
	#10 counter$count = 79953;
	#10 counter$count = 79954;
	#10 counter$count = 79955;
	#10 counter$count = 79956;
	#10 counter$count = 79957;
	#10 counter$count = 79958;
	#10 counter$count = 79959;
	#10 counter$count = 79960;
	#10 counter$count = 79961;
	#10 counter$count = 79962;
	#10 counter$count = 79963;
	#10 counter$count = 79964;
	#10 counter$count = 79965;
	#10 counter$count = 79966;
	#10 counter$count = 79967;
	#10 counter$count = 79968;
	#10 counter$count = 79969;
	#10 counter$count = 79970;
	#10 counter$count = 79971;
	#10 counter$count = 79972;
	#10 counter$count = 79973;
	#10 counter$count = 79974;
	#10 counter$count = 79975;
	#10 counter$count = 79976;
	#10 counter$count = 79977;
	#10 counter$count = 79978;
	#10 counter$count = 79979;
	#10 counter$count = 79980;
	#10 counter$count = 79981;
	#10 counter$count = 79982;
	#10 counter$count = 79983;
	#10 counter$count = 79984;
	#10 counter$count = 79985;
	#10 counter$count = 79986;
	#10 counter$count = 79987;
	#10 counter$count = 79988;
	#10 counter$count = 79989;
	#10 counter$count = 79990;
	#10 counter$count = 79991;
	#10 counter$count = 79992;
	#10 counter$count = 79993;
	#10 counter$count = 79994;
	#10 counter$count = 79995;
	#10 counter$count = 79996;
	#10 counter$count = 79997;
	#10 counter$count = 79998;
	#10 counter$count = 79999;
	#10 counter$count = 80000;
	#10 counter$count = 80001;
	#10 counter$count = 80002;
	#10 counter$count = 80003;
	#10 counter$count = 80004;
	#10 counter$count = 80005;
	#10 counter$count = 80006;
	#10 counter$count = 80007;
	#10 counter$count = 80008;
	#10 counter$count = 80009;
	#10 counter$count = 80010;
	#10 counter$count = 80011;
	#10 counter$count = 80012;
	#10 counter$count = 80013;
	#10 counter$count = 80014;
	#10 counter$count = 80015;
	#10 counter$count = 80016;
	#10 counter$count = 80017;
	#10 counter$count = 80018;
	#10 counter$count = 80019;
	#10 counter$count = 80020;
	#10 counter$count = 80021;
	#10 counter$count = 80022;
	#10 counter$count = 80023;
	#10 counter$count = 80024;
	#10 counter$count = 80025;
	#10 counter$count = 80026;
	#10 counter$count = 80027;
	#10 counter$count = 80028;
	#10 counter$count = 80029;
	#10 counter$count = 80030;
	#10 counter$count = 80031;
	#10 counter$count = 80032;
	#10 counter$count = 80033;
	#10 counter$count = 80034;
	#10 counter$count = 80035;
	#10 counter$count = 80036;
	#10 counter$count = 80037;
	#10 counter$count = 80038;
	#10 counter$count = 80039;
	#10 counter$count = 80040;
	#10 counter$count = 80041;
	#10 counter$count = 80042;
	#10 counter$count = 80043;
	#10 counter$count = 80044;
	#10 counter$count = 80045;
	#10 counter$count = 80046;
	#10 counter$count = 80047;
	#10 counter$count = 80048;
	#10 counter$count = 80049;
	#10 counter$count = 80050;
	#10 counter$count = 80051;
	#10 counter$count = 80052;
	#10 counter$count = 80053;
	#10 counter$count = 80054;
	#10 counter$count = 80055;
	#10 counter$count = 80056;
	#10 counter$count = 80057;
	#10 counter$count = 80058;
	#10 counter$count = 80059;
	#10 counter$count = 80060;
	#10 counter$count = 80061;
	#10 counter$count = 80062;
	#10 counter$count = 80063;
	#10 counter$count = 80064;
	#10 counter$count = 80065;
	#10 counter$count = 80066;
	#10 counter$count = 80067;
	#10 counter$count = 80068;
	#10 counter$count = 80069;
	#10 counter$count = 80070;
	#10 counter$count = 80071;
	#10 counter$count = 80072;
	#10 counter$count = 80073;
	#10 counter$count = 80074;
	#10 counter$count = 80075;
	#10 counter$count = 80076;
	#10 counter$count = 80077;
	#10 counter$count = 80078;
	#10 counter$count = 80079;
	#10 counter$count = 80080;
	#10 counter$count = 80081;
	#10 counter$count = 80082;
	#10 counter$count = 80083;
	#10 counter$count = 80084;
	#10 counter$count = 80085;
	#10 counter$count = 80086;
	#10 counter$count = 80087;
	#10 counter$count = 80088;
	#10 counter$count = 80089;
	#10 counter$count = 80090;
	#10 counter$count = 80091;
	#10 counter$count = 80092;
	#10 counter$count = 80093;
	#10 counter$count = 80094;
	#10 counter$count = 80095;
	#10 counter$count = 80096;
	#10 counter$count = 80097;
	#10 counter$count = 80098;
	#10 counter$count = 80099;
	#10 counter$count = 80100;
	#10 counter$count = 80101;
	#10 counter$count = 80102;
	#10 counter$count = 80103;
	#10 counter$count = 80104;
	#10 counter$count = 80105;
	#10 counter$count = 80106;
	#10 counter$count = 80107;
	#10 counter$count = 80108;
	#10 counter$count = 80109;
	#10 counter$count = 80110;
	#10 counter$count = 80111;
	#10 counter$count = 80112;
	#10 counter$count = 80113;
	#10 counter$count = 80114;
	#10 counter$count = 80115;
	#10 counter$count = 80116;
	#10 counter$count = 80117;
	#10 counter$count = 80118;
	#10 counter$count = 80119;
	#10 counter$count = 80120;
	#10 counter$count = 80121;
	#10 counter$count = 80122;
	#10 counter$count = 80123;
	#10 counter$count = 80124;
	#10 counter$count = 80125;
	#10 counter$count = 80126;
	#10 counter$count = 80127;
	#10 counter$count = 80128;
	#10 counter$count = 80129;
	#10 counter$count = 80130;
	#10 counter$count = 80131;
	#10 counter$count = 80132;
	#10 counter$count = 80133;
	#10 counter$count = 80134;
	#10 counter$count = 80135;
	#10 counter$count = 80136;
	#10 counter$count = 80137;
	#10 counter$count = 80138;
	#10 counter$count = 80139;
	#10 counter$count = 80140;
	#10 counter$count = 80141;
	#10 counter$count = 80142;
	#10 counter$count = 80143;
	#10 counter$count = 80144;
	#10 counter$count = 80145;
	#10 counter$count = 80146;
	#10 counter$count = 80147;
	#10 counter$count = 80148;
	#10 counter$count = 80149;
	#10 counter$count = 80150;
	#10 counter$count = 80151;
	#10 counter$count = 80152;
	#10 counter$count = 80153;
	#10 counter$count = 80154;
	#10 counter$count = 80155;
	#10 counter$count = 80156;
	#10 counter$count = 80157;
	#10 counter$count = 80158;
	#10 counter$count = 80159;
	#10 counter$count = 80160;
	#10 counter$count = 80161;
	#10 counter$count = 80162;
	#10 counter$count = 80163;
	#10 counter$count = 80164;
	#10 counter$count = 80165;
	#10 counter$count = 80166;
	#10 counter$count = 80167;
	#10 counter$count = 80168;
	#10 counter$count = 80169;
	#10 counter$count = 80170;
	#10 counter$count = 80171;
	#10 counter$count = 80172;
	#10 counter$count = 80173;
	#10 counter$count = 80174;
	#10 counter$count = 80175;
	#10 counter$count = 80176;
	#10 counter$count = 80177;
	#10 counter$count = 80178;
	#10 counter$count = 80179;
	#10 counter$count = 80180;
	#10 counter$count = 80181;
	#10 counter$count = 80182;
	#10 counter$count = 80183;
	#10 counter$count = 80184;
	#10 counter$count = 80185;
	#10 counter$count = 80186;
	#10 counter$count = 80187;
	#10 counter$count = 80188;
	#10 counter$count = 80189;
	#10 counter$count = 80190;
	#10 counter$count = 80191;
	#10 counter$count = 80192;
	#10 counter$count = 80193;
	#10 counter$count = 80194;
	#10 counter$count = 80195;
	#10 counter$count = 80196;
	#10 counter$count = 80197;
	#10 counter$count = 80198;
	#10 counter$count = 80199;
	#10 counter$count = 80200;
	#10 counter$count = 80201;
	#10 counter$count = 80202;
	#10 counter$count = 80203;
	#10 counter$count = 80204;
	#10 counter$count = 80205;
	#10 counter$count = 80206;
	#10 counter$count = 80207;
	#10 counter$count = 80208;
	#10 counter$count = 80209;
	#10 counter$count = 80210;
	#10 counter$count = 80211;
	#10 counter$count = 80212;
	#10 counter$count = 80213;
	#10 counter$count = 80214;
	#10 counter$count = 80215;
	#10 counter$count = 80216;
	#10 counter$count = 80217;
	#10 counter$count = 80218;
	#10 counter$count = 80219;
	#10 counter$count = 80220;
	#10 counter$count = 80221;
	#10 counter$count = 80222;
	#10 counter$count = 80223;
	#10 counter$count = 80224;
	#10 counter$count = 80225;
	#10 counter$count = 80226;
	#10 counter$count = 80227;
	#10 counter$count = 80228;
	#10 counter$count = 80229;
	#10 counter$count = 80230;
	#10 counter$count = 80231;
	#10 counter$count = 80232;
	#10 counter$count = 80233;
	#10 counter$count = 80234;
	#10 counter$count = 80235;
	#10 counter$count = 80236;
	#10 counter$count = 80237;
	#10 counter$count = 80238;
	#10 counter$count = 80239;
	#10 counter$count = 80240;
	#10 counter$count = 80241;
	#10 counter$count = 80242;
	#10 counter$count = 80243;
	#10 counter$count = 80244;
	#10 counter$count = 80245;
	#10 counter$count = 80246;
	#10 counter$count = 80247;
	#10 counter$count = 80248;
	#10 counter$count = 80249;
	#10 counter$count = 80250;
	#10 counter$count = 80251;
	#10 counter$count = 80252;
	#10 counter$count = 80253;
	#10 counter$count = 80254;
	#10 counter$count = 80255;
	#10 counter$count = 80256;
	#10 counter$count = 80257;
	#10 counter$count = 80258;
	#10 counter$count = 80259;
	#10 counter$count = 80260;
	#10 counter$count = 80261;
	#10 counter$count = 80262;
	#10 counter$count = 80263;
	#10 counter$count = 80264;
	#10 counter$count = 80265;
	#10 counter$count = 80266;
	#10 counter$count = 80267;
	#10 counter$count = 80268;
	#10 counter$count = 80269;
	#10 counter$count = 80270;
	#10 counter$count = 80271;
	#10 counter$count = 80272;
	#10 counter$count = 80273;
	#10 counter$count = 80274;
	#10 counter$count = 80275;
	#10 counter$count = 80276;
	#10 counter$count = 80277;
	#10 counter$count = 80278;
	#10 counter$count = 80279;
	#10 counter$count = 80280;
	#10 counter$count = 80281;
	#10 counter$count = 80282;
	#10 counter$count = 80283;
	#10 counter$count = 80284;
	#10 counter$count = 80285;
	#10 counter$count = 80286;
	#10 counter$count = 80287;
	#10 counter$count = 80288;
	#10 counter$count = 80289;
	#10 counter$count = 80290;
	#10 counter$count = 80291;
	#10 counter$count = 80292;
	#10 counter$count = 80293;
	#10 counter$count = 80294;
	#10 counter$count = 80295;
	#10 counter$count = 80296;
	#10 counter$count = 80297;
	#10 counter$count = 80298;
	#10 counter$count = 80299;
	#10 counter$count = 80300;
	#10 counter$count = 80301;
	#10 counter$count = 80302;
	#10 counter$count = 80303;
	#10 counter$count = 80304;
	#10 counter$count = 80305;
	#10 counter$count = 80306;
	#10 counter$count = 80307;
	#10 counter$count = 80308;
	#10 counter$count = 80309;
	#10 counter$count = 80310;
	#10 counter$count = 80311;
	#10 counter$count = 80312;
	#10 counter$count = 80313;
	#10 counter$count = 80314;
	#10 counter$count = 80315;
	#10 counter$count = 80316;
	#10 counter$count = 80317;
	#10 counter$count = 80318;
	#10 counter$count = 80319;
	#10 counter$count = 80320;
	#10 counter$count = 80321;
	#10 counter$count = 80322;
	#10 counter$count = 80323;
	#10 counter$count = 80324;
	#10 counter$count = 80325;
	#10 counter$count = 80326;
	#10 counter$count = 80327;
	#10 counter$count = 80328;
	#10 counter$count = 80329;
	#10 counter$count = 80330;
	#10 counter$count = 80331;
	#10 counter$count = 80332;
	#10 counter$count = 80333;
	#10 counter$count = 80334;
	#10 counter$count = 80335;
	#10 counter$count = 80336;
	#10 counter$count = 80337;
	#10 counter$count = 80338;
	#10 counter$count = 80339;
	#10 counter$count = 80340;
	#10 counter$count = 80341;
	#10 counter$count = 80342;
	#10 counter$count = 80343;
	#10 counter$count = 80344;
	#10 counter$count = 80345;
	#10 counter$count = 80346;
	#10 counter$count = 80347;
	#10 counter$count = 80348;
	#10 counter$count = 80349;
	#10 counter$count = 80350;
	#10 counter$count = 80351;
	#10 counter$count = 80352;
	#10 counter$count = 80353;
	#10 counter$count = 80354;
	#10 counter$count = 80355;
	#10 counter$count = 80356;
	#10 counter$count = 80357;
	#10 counter$count = 80358;
	#10 counter$count = 80359;
	#10 counter$count = 80360;
	#10 counter$count = 80361;
	#10 counter$count = 80362;
	#10 counter$count = 80363;
	#10 counter$count = 80364;
	#10 counter$count = 80365;
	#10 counter$count = 80366;
	#10 counter$count = 80367;
	#10 counter$count = 80368;
	#10 counter$count = 80369;
	#10 counter$count = 80370;
	#10 counter$count = 80371;
	#10 counter$count = 80372;
	#10 counter$count = 80373;
	#10 counter$count = 80374;
	#10 counter$count = 80375;
	#10 counter$count = 80376;
	#10 counter$count = 80377;
	#10 counter$count = 80378;
	#10 counter$count = 80379;
	#10 counter$count = 80380;
	#10 counter$count = 80381;
	#10 counter$count = 80382;
	#10 counter$count = 80383;
	#10 counter$count = 80384;
	#10 counter$count = 80385;
	#10 counter$count = 80386;
	#10 counter$count = 80387;
	#10 counter$count = 80388;
	#10 counter$count = 80389;
	#10 counter$count = 80390;
	#10 counter$count = 80391;
	#10 counter$count = 80392;
	#10 counter$count = 80393;
	#10 counter$count = 80394;
	#10 counter$count = 80395;
	#10 counter$count = 80396;
	#10 counter$count = 80397;
	#10 counter$count = 80398;
	#10 counter$count = 80399;
	#10 counter$count = 80400;
	#10 counter$count = 80401;
	#10 counter$count = 80402;
	#10 counter$count = 80403;
	#10 counter$count = 80404;
	#10 counter$count = 80405;
	#10 counter$count = 80406;
	#10 counter$count = 80407;
	#10 counter$count = 80408;
	#10 counter$count = 80409;
	#10 counter$count = 80410;
	#10 counter$count = 80411;
	#10 counter$count = 80412;
	#10 counter$count = 80413;
	#10 counter$count = 80414;
	#10 counter$count = 80415;
	#10 counter$count = 80416;
	#10 counter$count = 80417;
	#10 counter$count = 80418;
	#10 counter$count = 80419;
	#10 counter$count = 80420;
	#10 counter$count = 80421;
	#10 counter$count = 80422;
	#10 counter$count = 80423;
	#10 counter$count = 80424;
	#10 counter$count = 80425;
	#10 counter$count = 80426;
	#10 counter$count = 80427;
	#10 counter$count = 80428;
	#10 counter$count = 80429;
	#10 counter$count = 80430;
	#10 counter$count = 80431;
	#10 counter$count = 80432;
	#10 counter$count = 80433;
	#10 counter$count = 80434;
	#10 counter$count = 80435;
	#10 counter$count = 80436;
	#10 counter$count = 80437;
	#10 counter$count = 80438;
	#10 counter$count = 80439;
	#10 counter$count = 80440;
	#10 counter$count = 80441;
	#10 counter$count = 80442;
	#10 counter$count = 80443;
	#10 counter$count = 80444;
	#10 counter$count = 80445;
	#10 counter$count = 80446;
	#10 counter$count = 80447;
	#10 counter$count = 80448;
	#10 counter$count = 80449;
	#10 counter$count = 80450;
	#10 counter$count = 80451;
	#10 counter$count = 80452;
	#10 counter$count = 80453;
	#10 counter$count = 80454;
	#10 counter$count = 80455;
	#10 counter$count = 80456;
	#10 counter$count = 80457;
	#10 counter$count = 80458;
	#10 counter$count = 80459;
	#10 counter$count = 80460;
	#10 counter$count = 80461;
	#10 counter$count = 80462;
	#10 counter$count = 80463;
	#10 counter$count = 80464;
	#10 counter$count = 80465;
	#10 counter$count = 80466;
	#10 counter$count = 80467;
	#10 counter$count = 80468;
	#10 counter$count = 80469;
	#10 counter$count = 80470;
	#10 counter$count = 80471;
	#10 counter$count = 80472;
	#10 counter$count = 80473;
	#10 counter$count = 80474;
	#10 counter$count = 80475;
	#10 counter$count = 80476;
	#10 counter$count = 80477;
	#10 counter$count = 80478;
	#10 counter$count = 80479;
	#10 counter$count = 80480;
	#10 counter$count = 80481;
	#10 counter$count = 80482;
	#10 counter$count = 80483;
	#10 counter$count = 80484;
	#10 counter$count = 80485;
	#10 counter$count = 80486;
	#10 counter$count = 80487;
	#10 counter$count = 80488;
	#10 counter$count = 80489;
	#10 counter$count = 80490;
	#10 counter$count = 80491;
	#10 counter$count = 80492;
	#10 counter$count = 80493;
	#10 counter$count = 80494;
	#10 counter$count = 80495;
	#10 counter$count = 80496;
	#10 counter$count = 80497;
	#10 counter$count = 80498;
	#10 counter$count = 80499;
	#10 counter$count = 80500;
	#10 counter$count = 80501;
	#10 counter$count = 80502;
	#10 counter$count = 80503;
	#10 counter$count = 80504;
	#10 counter$count = 80505;
	#10 counter$count = 80506;
	#10 counter$count = 80507;
	#10 counter$count = 80508;
	#10 counter$count = 80509;
	#10 counter$count = 80510;
	#10 counter$count = 80511;
	#10 counter$count = 80512;
	#10 counter$count = 80513;
	#10 counter$count = 80514;
	#10 counter$count = 80515;
	#10 counter$count = 80516;
	#10 counter$count = 80517;
	#10 counter$count = 80518;
	#10 counter$count = 80519;
	#10 counter$count = 80520;
	#10 counter$count = 80521;
	#10 counter$count = 80522;
	#10 counter$count = 80523;
	#10 counter$count = 80524;
	#10 counter$count = 80525;
	#10 counter$count = 80526;
	#10 counter$count = 80527;
	#10 counter$count = 80528;
	#10 counter$count = 80529;
	#10 counter$count = 80530;
	#10 counter$count = 80531;
	#10 counter$count = 80532;
	#10 counter$count = 80533;
	#10 counter$count = 80534;
	#10 counter$count = 80535;
	#10 counter$count = 80536;
	#10 counter$count = 80537;
	#10 counter$count = 80538;
	#10 counter$count = 80539;
	#10 counter$count = 80540;
	#10 counter$count = 80541;
	#10 counter$count = 80542;
	#10 counter$count = 80543;
	#10 counter$count = 80544;
	#10 counter$count = 80545;
	#10 counter$count = 80546;
	#10 counter$count = 80547;
	#10 counter$count = 80548;
	#10 counter$count = 80549;
	#10 counter$count = 80550;
	#10 counter$count = 80551;
	#10 counter$count = 80552;
	#10 counter$count = 80553;
	#10 counter$count = 80554;
	#10 counter$count = 80555;
	#10 counter$count = 80556;
	#10 counter$count = 80557;
	#10 counter$count = 80558;
	#10 counter$count = 80559;
	#10 counter$count = 80560;
	#10 counter$count = 80561;
	#10 counter$count = 80562;
	#10 counter$count = 80563;
	#10 counter$count = 80564;
	#10 counter$count = 80565;
	#10 counter$count = 80566;
	#10 counter$count = 80567;
	#10 counter$count = 80568;
	#10 counter$count = 80569;
	#10 counter$count = 80570;
	#10 counter$count = 80571;
	#10 counter$count = 80572;
	#10 counter$count = 80573;
	#10 counter$count = 80574;
	#10 counter$count = 80575;
	#10 counter$count = 80576;
	#10 counter$count = 80577;
	#10 counter$count = 80578;
	#10 counter$count = 80579;
	#10 counter$count = 80580;
	#10 counter$count = 80581;
	#10 counter$count = 80582;
	#10 counter$count = 80583;
	#10 counter$count = 80584;
	#10 counter$count = 80585;
	#10 counter$count = 80586;
	#10 counter$count = 80587;
	#10 counter$count = 80588;
	#10 counter$count = 80589;
	#10 counter$count = 80590;
	#10 counter$count = 80591;
	#10 counter$count = 80592;
	#10 counter$count = 80593;
	#10 counter$count = 80594;
	#10 counter$count = 80595;
	#10 counter$count = 80596;
	#10 counter$count = 80597;
	#10 counter$count = 80598;
	#10 counter$count = 80599;
	#10 counter$count = 80600;
	#10 counter$count = 80601;
	#10 counter$count = 80602;
	#10 counter$count = 80603;
	#10 counter$count = 80604;
	#10 counter$count = 80605;
	#10 counter$count = 80606;
	#10 counter$count = 80607;
	#10 counter$count = 80608;
	#10 counter$count = 80609;
	#10 counter$count = 80610;
	#10 counter$count = 80611;
	#10 counter$count = 80612;
	#10 counter$count = 80613;
	#10 counter$count = 80614;
	#10 counter$count = 80615;
	#10 counter$count = 80616;
	#10 counter$count = 80617;
	#10 counter$count = 80618;
	#10 counter$count = 80619;
	#10 counter$count = 80620;
	#10 counter$count = 80621;
	#10 counter$count = 80622;
	#10 counter$count = 80623;
	#10 counter$count = 80624;
	#10 counter$count = 80625;
	#10 counter$count = 80626;
	#10 counter$count = 80627;
	#10 counter$count = 80628;
	#10 counter$count = 80629;
	#10 counter$count = 80630;
	#10 counter$count = 80631;
	#10 counter$count = 80632;
	#10 counter$count = 80633;
	#10 counter$count = 80634;
	#10 counter$count = 80635;
	#10 counter$count = 80636;
	#10 counter$count = 80637;
	#10 counter$count = 80638;
	#10 counter$count = 80639;
	#10 counter$count = 80640;
	#10 counter$count = 80641;
	#10 counter$count = 80642;
	#10 counter$count = 80643;
	#10 counter$count = 80644;
	#10 counter$count = 80645;
	#10 counter$count = 80646;
	#10 counter$count = 80647;
	#10 counter$count = 80648;
	#10 counter$count = 80649;
	#10 counter$count = 80650;
	#10 counter$count = 80651;
	#10 counter$count = 80652;
	#10 counter$count = 80653;
	#10 counter$count = 80654;
	#10 counter$count = 80655;
	#10 counter$count = 80656;
	#10 counter$count = 80657;
	#10 counter$count = 80658;
	#10 counter$count = 80659;
	#10 counter$count = 80660;
	#10 counter$count = 80661;
	#10 counter$count = 80662;
	#10 counter$count = 80663;
	#10 counter$count = 80664;
	#10 counter$count = 80665;
	#10 counter$count = 80666;
	#10 counter$count = 80667;
	#10 counter$count = 80668;
	#10 counter$count = 80669;
	#10 counter$count = 80670;
	#10 counter$count = 80671;
	#10 counter$count = 80672;
	#10 counter$count = 80673;
	#10 counter$count = 80674;
	#10 counter$count = 80675;
	#10 counter$count = 80676;
	#10 counter$count = 80677;
	#10 counter$count = 80678;
	#10 counter$count = 80679;
	#10 counter$count = 80680;
	#10 counter$count = 80681;
	#10 counter$count = 80682;
	#10 counter$count = 80683;
	#10 counter$count = 80684;
	#10 counter$count = 80685;
	#10 counter$count = 80686;
	#10 counter$count = 80687;
	#10 counter$count = 80688;
	#10 counter$count = 80689;
	#10 counter$count = 80690;
	#10 counter$count = 80691;
	#10 counter$count = 80692;
	#10 counter$count = 80693;
	#10 counter$count = 80694;
	#10 counter$count = 80695;
	#10 counter$count = 80696;
	#10 counter$count = 80697;
	#10 counter$count = 80698;
	#10 counter$count = 80699;
	#10 counter$count = 80700;
	#10 counter$count = 80701;
	#10 counter$count = 80702;
	#10 counter$count = 80703;
	#10 counter$count = 80704;
	#10 counter$count = 80705;
	#10 counter$count = 80706;
	#10 counter$count = 80707;
	#10 counter$count = 80708;
	#10 counter$count = 80709;
	#10 counter$count = 80710;
	#10 counter$count = 80711;
	#10 counter$count = 80712;
	#10 counter$count = 80713;
	#10 counter$count = 80714;
	#10 counter$count = 80715;
	#10 counter$count = 80716;
	#10 counter$count = 80717;
	#10 counter$count = 80718;
	#10 counter$count = 80719;
	#10 counter$count = 80720;
	#10 counter$count = 80721;
	#10 counter$count = 80722;
	#10 counter$count = 80723;
	#10 counter$count = 80724;
	#10 counter$count = 80725;
	#10 counter$count = 80726;
	#10 counter$count = 80727;
	#10 counter$count = 80728;
	#10 counter$count = 80729;
	#10 counter$count = 80730;
	#10 counter$count = 80731;
	#10 counter$count = 80732;
	#10 counter$count = 80733;
	#10 counter$count = 80734;
	#10 counter$count = 80735;
	#10 counter$count = 80736;
	#10 counter$count = 80737;
	#10 counter$count = 80738;
	#10 counter$count = 80739;
	#10 counter$count = 80740;
	#10 counter$count = 80741;
	#10 counter$count = 80742;
	#10 counter$count = 80743;
	#10 counter$count = 80744;
	#10 counter$count = 80745;
	#10 counter$count = 80746;
	#10 counter$count = 80747;
	#10 counter$count = 80748;
	#10 counter$count = 80749;
	#10 counter$count = 80750;
	#10 counter$count = 80751;
	#10 counter$count = 80752;
	#10 counter$count = 80753;
	#10 counter$count = 80754;
	#10 counter$count = 80755;
	#10 counter$count = 80756;
	#10 counter$count = 80757;
	#10 counter$count = 80758;
	#10 counter$count = 80759;
	#10 counter$count = 80760;
	#10 counter$count = 80761;
	#10 counter$count = 80762;
	#10 counter$count = 80763;
	#10 counter$count = 80764;
	#10 counter$count = 80765;
	#10 counter$count = 80766;
	#10 counter$count = 80767;
	#10 counter$count = 80768;
	#10 counter$count = 80769;
	#10 counter$count = 80770;
	#10 counter$count = 80771;
	#10 counter$count = 80772;
	#10 counter$count = 80773;
	#10 counter$count = 80774;
	#10 counter$count = 80775;
	#10 counter$count = 80776;
	#10 counter$count = 80777;
	#10 counter$count = 80778;
	#10 counter$count = 80779;
	#10 counter$count = 80780;
	#10 counter$count = 80781;
	#10 counter$count = 80782;
	#10 counter$count = 80783;
	#10 counter$count = 80784;
	#10 counter$count = 80785;
	#10 counter$count = 80786;
	#10 counter$count = 80787;
	#10 counter$count = 80788;
	#10 counter$count = 80789;
	#10 counter$count = 80790;
	#10 counter$count = 80791;
	#10 counter$count = 80792;
	#10 counter$count = 80793;
	#10 counter$count = 80794;
	#10 counter$count = 80795;
	#10 counter$count = 80796;
	#10 counter$count = 80797;
	#10 counter$count = 80798;
	#10 counter$count = 80799;
	#10 counter$count = 80800;
	#10 counter$count = 80801;
	#10 counter$count = 80802;
	#10 counter$count = 80803;
	#10 counter$count = 80804;
	#10 counter$count = 80805;
	#10 counter$count = 80806;
	#10 counter$count = 80807;
	#10 counter$count = 80808;
	#10 counter$count = 80809;
	#10 counter$count = 80810;
	#10 counter$count = 80811;
	#10 counter$count = 80812;
	#10 counter$count = 80813;
	#10 counter$count = 80814;
	#10 counter$count = 80815;
	#10 counter$count = 80816;
	#10 counter$count = 80817;
	#10 counter$count = 80818;
	#10 counter$count = 80819;
	#10 counter$count = 80820;
	#10 counter$count = 80821;
	#10 counter$count = 80822;
	#10 counter$count = 80823;
	#10 counter$count = 80824;
	#10 counter$count = 80825;
	#10 counter$count = 80826;
	#10 counter$count = 80827;
	#10 counter$count = 80828;
	#10 counter$count = 80829;
	#10 counter$count = 80830;
	#10 counter$count = 80831;
	#10 counter$count = 80832;
	#10 counter$count = 80833;
	#10 counter$count = 80834;
	#10 counter$count = 80835;
	#10 counter$count = 80836;
	#10 counter$count = 80837;
	#10 counter$count = 80838;
	#10 counter$count = 80839;
	#10 counter$count = 80840;
	#10 counter$count = 80841;
	#10 counter$count = 80842;
	#10 counter$count = 80843;
	#10 counter$count = 80844;
	#10 counter$count = 80845;
	#10 counter$count = 80846;
	#10 counter$count = 80847;
	#10 counter$count = 80848;
	#10 counter$count = 80849;
	#10 counter$count = 80850;
	#10 counter$count = 80851;
	#10 counter$count = 80852;
	#10 counter$count = 80853;
	#10 counter$count = 80854;
	#10 counter$count = 80855;
	#10 counter$count = 80856;
	#10 counter$count = 80857;
	#10 counter$count = 80858;
	#10 counter$count = 80859;
	#10 counter$count = 80860;
	#10 counter$count = 80861;
	#10 counter$count = 80862;
	#10 counter$count = 80863;
	#10 counter$count = 80864;
	#10 counter$count = 80865;
	#10 counter$count = 80866;
	#10 counter$count = 80867;
	#10 counter$count = 80868;
	#10 counter$count = 80869;
	#10 counter$count = 80870;
	#10 counter$count = 80871;
	#10 counter$count = 80872;
	#10 counter$count = 80873;
	#10 counter$count = 80874;
	#10 counter$count = 80875;
	#10 counter$count = 80876;
	#10 counter$count = 80877;
	#10 counter$count = 80878;
	#10 counter$count = 80879;
	#10 counter$count = 80880;
	#10 counter$count = 80881;
	#10 counter$count = 80882;
	#10 counter$count = 80883;
	#10 counter$count = 80884;
	#10 counter$count = 80885;
	#10 counter$count = 80886;
	#10 counter$count = 80887;
	#10 counter$count = 80888;
	#10 counter$count = 80889;
	#10 counter$count = 80890;
	#10 counter$count = 80891;
	#10 counter$count = 80892;
	#10 counter$count = 80893;
	#10 counter$count = 80894;
	#10 counter$count = 80895;
	#10 counter$count = 80896;
	#10 counter$count = 80897;
	#10 counter$count = 80898;
	#10 counter$count = 80899;
	#10 counter$count = 80900;
	#10 counter$count = 80901;
	#10 counter$count = 80902;
	#10 counter$count = 80903;
	#10 counter$count = 80904;
	#10 counter$count = 80905;
	#10 counter$count = 80906;
	#10 counter$count = 80907;
	#10 counter$count = 80908;
	#10 counter$count = 80909;
	#10 counter$count = 80910;
	#10 counter$count = 80911;
	#10 counter$count = 80912;
	#10 counter$count = 80913;
	#10 counter$count = 80914;
	#10 counter$count = 80915;
	#10 counter$count = 80916;
	#10 counter$count = 80917;
	#10 counter$count = 80918;
	#10 counter$count = 80919;
	#10 counter$count = 80920;
	#10 counter$count = 80921;
	#10 counter$count = 80922;
	#10 counter$count = 80923;
	#10 counter$count = 80924;
	#10 counter$count = 80925;
	#10 counter$count = 80926;
	#10 counter$count = 80927;
	#10 counter$count = 80928;
	#10 counter$count = 80929;
	#10 counter$count = 80930;
	#10 counter$count = 80931;
	#10 counter$count = 80932;
	#10 counter$count = 80933;
	#10 counter$count = 80934;
	#10 counter$count = 80935;
	#10 counter$count = 80936;
	#10 counter$count = 80937;
	#10 counter$count = 80938;
	#10 counter$count = 80939;
	#10 counter$count = 80940;
	#10 counter$count = 80941;
	#10 counter$count = 80942;
	#10 counter$count = 80943;
	#10 counter$count = 80944;
	#10 counter$count = 80945;
	#10 counter$count = 80946;
	#10 counter$count = 80947;
	#10 counter$count = 80948;
	#10 counter$count = 80949;
	#10 counter$count = 80950;
	#10 counter$count = 80951;
	#10 counter$count = 80952;
	#10 counter$count = 80953;
	#10 counter$count = 80954;
	#10 counter$count = 80955;
	#10 counter$count = 80956;
	#10 counter$count = 80957;
	#10 counter$count = 80958;
	#10 counter$count = 80959;
	#10 counter$count = 80960;
	#10 counter$count = 80961;
	#10 counter$count = 80962;
	#10 counter$count = 80963;
	#10 counter$count = 80964;
	#10 counter$count = 80965;
	#10 counter$count = 80966;
	#10 counter$count = 80967;
	#10 counter$count = 80968;
	#10 counter$count = 80969;
	#10 counter$count = 80970;
	#10 counter$count = 80971;
	#10 counter$count = 80972;
	#10 counter$count = 80973;
	#10 counter$count = 80974;
	#10 counter$count = 80975;
	#10 counter$count = 80976;
	#10 counter$count = 80977;
	#10 counter$count = 80978;
	#10 counter$count = 80979;
	#10 counter$count = 80980;
	#10 counter$count = 80981;
	#10 counter$count = 80982;
	#10 counter$count = 80983;
	#10 counter$count = 80984;
	#10 counter$count = 80985;
	#10 counter$count = 80986;
	#10 counter$count = 80987;
	#10 counter$count = 80988;
	#10 counter$count = 80989;
	#10 counter$count = 80990;
	#10 counter$count = 80991;
	#10 counter$count = 80992;
	#10 counter$count = 80993;
	#10 counter$count = 80994;
	#10 counter$count = 80995;
	#10 counter$count = 80996;
	#10 counter$count = 80997;
	#10 counter$count = 80998;
	#10 counter$count = 80999;
	#10 counter$count = 81000;
	#10 counter$count = 81001;
	#10 counter$count = 81002;
	#10 counter$count = 81003;
	#10 counter$count = 81004;
	#10 counter$count = 81005;
	#10 counter$count = 81006;
	#10 counter$count = 81007;
	#10 counter$count = 81008;
	#10 counter$count = 81009;
	#10 counter$count = 81010;
	#10 counter$count = 81011;
	#10 counter$count = 81012;
	#10 counter$count = 81013;
	#10 counter$count = 81014;
	#10 counter$count = 81015;
	#10 counter$count = 81016;
	#10 counter$count = 81017;
	#10 counter$count = 81018;
	#10 counter$count = 81019;
	#10 counter$count = 81020;
	#10 counter$count = 81021;
	#10 counter$count = 81022;
	#10 counter$count = 81023;
	#10 counter$count = 81024;
	#10 counter$count = 81025;
	#10 counter$count = 81026;
	#10 counter$count = 81027;
	#10 counter$count = 81028;
	#10 counter$count = 81029;
	#10 counter$count = 81030;
	#10 counter$count = 81031;
	#10 counter$count = 81032;
	#10 counter$count = 81033;
	#10 counter$count = 81034;
	#10 counter$count = 81035;
	#10 counter$count = 81036;
	#10 counter$count = 81037;
	#10 counter$count = 81038;
	#10 counter$count = 81039;
	#10 counter$count = 81040;
	#10 counter$count = 81041;
	#10 counter$count = 81042;
	#10 counter$count = 81043;
	#10 counter$count = 81044;
	#10 counter$count = 81045;
	#10 counter$count = 81046;
	#10 counter$count = 81047;
	#10 counter$count = 81048;
	#10 counter$count = 81049;
	#10 counter$count = 81050;
	#10 counter$count = 81051;
	#10 counter$count = 81052;
	#10 counter$count = 81053;
	#10 counter$count = 81054;
	#10 counter$count = 81055;
	#10 counter$count = 81056;
	#10 counter$count = 81057;
	#10 counter$count = 81058;
	#10 counter$count = 81059;
	#10 counter$count = 81060;
	#10 counter$count = 81061;
	#10 counter$count = 81062;
	#10 counter$count = 81063;
	#10 counter$count = 81064;
	#10 counter$count = 81065;
	#10 counter$count = 81066;
	#10 counter$count = 81067;
	#10 counter$count = 81068;
	#10 counter$count = 81069;
	#10 counter$count = 81070;
	#10 counter$count = 81071;
	#10 counter$count = 81072;
	#10 counter$count = 81073;
	#10 counter$count = 81074;
	#10 counter$count = 81075;
	#10 counter$count = 81076;
	#10 counter$count = 81077;
	#10 counter$count = 81078;
	#10 counter$count = 81079;
	#10 counter$count = 81080;
	#10 counter$count = 81081;
	#10 counter$count = 81082;
	#10 counter$count = 81083;
	#10 counter$count = 81084;
	#10 counter$count = 81085;
	#10 counter$count = 81086;
	#10 counter$count = 81087;
	#10 counter$count = 81088;
	#10 counter$count = 81089;
	#10 counter$count = 81090;
	#10 counter$count = 81091;
	#10 counter$count = 81092;
	#10 counter$count = 81093;
	#10 counter$count = 81094;
	#10 counter$count = 81095;
	#10 counter$count = 81096;
	#10 counter$count = 81097;
	#10 counter$count = 81098;
	#10 counter$count = 81099;
	#10 counter$count = 81100;
	#10 counter$count = 81101;
	#10 counter$count = 81102;
	#10 counter$count = 81103;
	#10 counter$count = 81104;
	#10 counter$count = 81105;
	#10 counter$count = 81106;
	#10 counter$count = 81107;
	#10 counter$count = 81108;
	#10 counter$count = 81109;
	#10 counter$count = 81110;
	#10 counter$count = 81111;
	#10 counter$count = 81112;
	#10 counter$count = 81113;
	#10 counter$count = 81114;
	#10 counter$count = 81115;
	#10 counter$count = 81116;
	#10 counter$count = 81117;
	#10 counter$count = 81118;
	#10 counter$count = 81119;
	#10 counter$count = 81120;
	#10 counter$count = 81121;
	#10 counter$count = 81122;
	#10 counter$count = 81123;
	#10 counter$count = 81124;
	#10 counter$count = 81125;
	#10 counter$count = 81126;
	#10 counter$count = 81127;
	#10 counter$count = 81128;
	#10 counter$count = 81129;
	#10 counter$count = 81130;
	#10 counter$count = 81131;
	#10 counter$count = 81132;
	#10 counter$count = 81133;
	#10 counter$count = 81134;
	#10 counter$count = 81135;
	#10 counter$count = 81136;
	#10 counter$count = 81137;
	#10 counter$count = 81138;
	#10 counter$count = 81139;
	#10 counter$count = 81140;
	#10 counter$count = 81141;
	#10 counter$count = 81142;
	#10 counter$count = 81143;
	#10 counter$count = 81144;
	#10 counter$count = 81145;
	#10 counter$count = 81146;
	#10 counter$count = 81147;
	#10 counter$count = 81148;
	#10 counter$count = 81149;
	#10 counter$count = 81150;
	#10 counter$count = 81151;
	#10 counter$count = 81152;
	#10 counter$count = 81153;
	#10 counter$count = 81154;
	#10 counter$count = 81155;
	#10 counter$count = 81156;
	#10 counter$count = 81157;
	#10 counter$count = 81158;
	#10 counter$count = 81159;
	#10 counter$count = 81160;
	#10 counter$count = 81161;
	#10 counter$count = 81162;
	#10 counter$count = 81163;
	#10 counter$count = 81164;
	#10 counter$count = 81165;
	#10 counter$count = 81166;
	#10 counter$count = 81167;
	#10 counter$count = 81168;
	#10 counter$count = 81169;
	#10 counter$count = 81170;
	#10 counter$count = 81171;
	#10 counter$count = 81172;
	#10 counter$count = 81173;
	#10 counter$count = 81174;
	#10 counter$count = 81175;
	#10 counter$count = 81176;
	#10 counter$count = 81177;
	#10 counter$count = 81178;
	#10 counter$count = 81179;
	#10 counter$count = 81180;
	#10 counter$count = 81181;
	#10 counter$count = 81182;
	#10 counter$count = 81183;
	#10 counter$count = 81184;
	#10 counter$count = 81185;
	#10 counter$count = 81186;
	#10 counter$count = 81187;
	#10 counter$count = 81188;
	#10 counter$count = 81189;
	#10 counter$count = 81190;
	#10 counter$count = 81191;
	#10 counter$count = 81192;
	#10 counter$count = 81193;
	#10 counter$count = 81194;
	#10 counter$count = 81195;
	#10 counter$count = 81196;
	#10 counter$count = 81197;
	#10 counter$count = 81198;
	#10 counter$count = 81199;
	#10 counter$count = 81200;
	#10 counter$count = 81201;
	#10 counter$count = 81202;
	#10 counter$count = 81203;
	#10 counter$count = 81204;
	#10 counter$count = 81205;
	#10 counter$count = 81206;
	#10 counter$count = 81207;
	#10 counter$count = 81208;
	#10 counter$count = 81209;
	#10 counter$count = 81210;
	#10 counter$count = 81211;
	#10 counter$count = 81212;
	#10 counter$count = 81213;
	#10 counter$count = 81214;
	#10 counter$count = 81215;
	#10 counter$count = 81216;
	#10 counter$count = 81217;
	#10 counter$count = 81218;
	#10 counter$count = 81219;
	#10 counter$count = 81220;
	#10 counter$count = 81221;
	#10 counter$count = 81222;
	#10 counter$count = 81223;
	#10 counter$count = 81224;
	#10 counter$count = 81225;
	#10 counter$count = 81226;
	#10 counter$count = 81227;
	#10 counter$count = 81228;
	#10 counter$count = 81229;
	#10 counter$count = 81230;
	#10 counter$count = 81231;
	#10 counter$count = 81232;
	#10 counter$count = 81233;
	#10 counter$count = 81234;
	#10 counter$count = 81235;
	#10 counter$count = 81236;
	#10 counter$count = 81237;
	#10 counter$count = 81238;
	#10 counter$count = 81239;
	#10 counter$count = 81240;
	#10 counter$count = 81241;
	#10 counter$count = 81242;
	#10 counter$count = 81243;
	#10 counter$count = 81244;
	#10 counter$count = 81245;
	#10 counter$count = 81246;
	#10 counter$count = 81247;
	#10 counter$count = 81248;
	#10 counter$count = 81249;
	#10 counter$count = 81250;
	#10 counter$count = 81251;
	#10 counter$count = 81252;
	#10 counter$count = 81253;
	#10 counter$count = 81254;
	#10 counter$count = 81255;
	#10 counter$count = 81256;
	#10 counter$count = 81257;
	#10 counter$count = 81258;
	#10 counter$count = 81259;
	#10 counter$count = 81260;
	#10 counter$count = 81261;
	#10 counter$count = 81262;
	#10 counter$count = 81263;
	#10 counter$count = 81264;
	#10 counter$count = 81265;
	#10 counter$count = 81266;
	#10 counter$count = 81267;
	#10 counter$count = 81268;
	#10 counter$count = 81269;
	#10 counter$count = 81270;
	#10 counter$count = 81271;
	#10 counter$count = 81272;
	#10 counter$count = 81273;
	#10 counter$count = 81274;
	#10 counter$count = 81275;
	#10 counter$count = 81276;
	#10 counter$count = 81277;
	#10 counter$count = 81278;
	#10 counter$count = 81279;
	#10 counter$count = 81280;
	#10 counter$count = 81281;
	#10 counter$count = 81282;
	#10 counter$count = 81283;
	#10 counter$count = 81284;
	#10 counter$count = 81285;
	#10 counter$count = 81286;
	#10 counter$count = 81287;
	#10 counter$count = 81288;
	#10 counter$count = 81289;
	#10 counter$count = 81290;
	#10 counter$count = 81291;
	#10 counter$count = 81292;
	#10 counter$count = 81293;
	#10 counter$count = 81294;
	#10 counter$count = 81295;
	#10 counter$count = 81296;
	#10 counter$count = 81297;
	#10 counter$count = 81298;
	#10 counter$count = 81299;
	#10 counter$count = 81300;
	#10 counter$count = 81301;
	#10 counter$count = 81302;
	#10 counter$count = 81303;
	#10 counter$count = 81304;
	#10 counter$count = 81305;
	#10 counter$count = 81306;
	#10 counter$count = 81307;
	#10 counter$count = 81308;
	#10 counter$count = 81309;
	#10 counter$count = 81310;
	#10 counter$count = 81311;
	#10 counter$count = 81312;
	#10 counter$count = 81313;
	#10 counter$count = 81314;
	#10 counter$count = 81315;
	#10 counter$count = 81316;
	#10 counter$count = 81317;
	#10 counter$count = 81318;
	#10 counter$count = 81319;
	#10 counter$count = 81320;
	#10 counter$count = 81321;
	#10 counter$count = 81322;
	#10 counter$count = 81323;
	#10 counter$count = 81324;
	#10 counter$count = 81325;
	#10 counter$count = 81326;
	#10 counter$count = 81327;
	#10 counter$count = 81328;
	#10 counter$count = 81329;
	#10 counter$count = 81330;
	#10 counter$count = 81331;
	#10 counter$count = 81332;
	#10 counter$count = 81333;
	#10 counter$count = 81334;
	#10 counter$count = 81335;
	#10 counter$count = 81336;
	#10 counter$count = 81337;
	#10 counter$count = 81338;
	#10 counter$count = 81339;
	#10 counter$count = 81340;
	#10 counter$count = 81341;
	#10 counter$count = 81342;
	#10 counter$count = 81343;
	#10 counter$count = 81344;
	#10 counter$count = 81345;
	#10 counter$count = 81346;
	#10 counter$count = 81347;
	#10 counter$count = 81348;
	#10 counter$count = 81349;
	#10 counter$count = 81350;
	#10 counter$count = 81351;
	#10 counter$count = 81352;
	#10 counter$count = 81353;
	#10 counter$count = 81354;
	#10 counter$count = 81355;
	#10 counter$count = 81356;
	#10 counter$count = 81357;
	#10 counter$count = 81358;
	#10 counter$count = 81359;
	#10 counter$count = 81360;
	#10 counter$count = 81361;
	#10 counter$count = 81362;
	#10 counter$count = 81363;
	#10 counter$count = 81364;
	#10 counter$count = 81365;
	#10 counter$count = 81366;
	#10 counter$count = 81367;
	#10 counter$count = 81368;
	#10 counter$count = 81369;
	#10 counter$count = 81370;
	#10 counter$count = 81371;
	#10 counter$count = 81372;
	#10 counter$count = 81373;
	#10 counter$count = 81374;
	#10 counter$count = 81375;
	#10 counter$count = 81376;
	#10 counter$count = 81377;
	#10 counter$count = 81378;
	#10 counter$count = 81379;
	#10 counter$count = 81380;
	#10 counter$count = 81381;
	#10 counter$count = 81382;
	#10 counter$count = 81383;
	#10 counter$count = 81384;
	#10 counter$count = 81385;
	#10 counter$count = 81386;
	#10 counter$count = 81387;
	#10 counter$count = 81388;
	#10 counter$count = 81389;
	#10 counter$count = 81390;
	#10 counter$count = 81391;
	#10 counter$count = 81392;
	#10 counter$count = 81393;
	#10 counter$count = 81394;
	#10 counter$count = 81395;
	#10 counter$count = 81396;
	#10 counter$count = 81397;
	#10 counter$count = 81398;
	#10 counter$count = 81399;
	#10 counter$count = 81400;
	#10 counter$count = 81401;
	#10 counter$count = 81402;
	#10 counter$count = 81403;
	#10 counter$count = 81404;
	#10 counter$count = 81405;
	#10 counter$count = 81406;
	#10 counter$count = 81407;
	#10 counter$count = 81408;
	#10 counter$count = 81409;
	#10 counter$count = 81410;
	#10 counter$count = 81411;
	#10 counter$count = 81412;
	#10 counter$count = 81413;
	#10 counter$count = 81414;
	#10 counter$count = 81415;
	#10 counter$count = 81416;
	#10 counter$count = 81417;
	#10 counter$count = 81418;
	#10 counter$count = 81419;
	#10 counter$count = 81420;
	#10 counter$count = 81421;
	#10 counter$count = 81422;
	#10 counter$count = 81423;
	#10 counter$count = 81424;
	#10 counter$count = 81425;
	#10 counter$count = 81426;
	#10 counter$count = 81427;
	#10 counter$count = 81428;
	#10 counter$count = 81429;
	#10 counter$count = 81430;
	#10 counter$count = 81431;
	#10 counter$count = 81432;
	#10 counter$count = 81433;
	#10 counter$count = 81434;
	#10 counter$count = 81435;
	#10 counter$count = 81436;
	#10 counter$count = 81437;
	#10 counter$count = 81438;
	#10 counter$count = 81439;
	#10 counter$count = 81440;
	#10 counter$count = 81441;
	#10 counter$count = 81442;
	#10 counter$count = 81443;
	#10 counter$count = 81444;
	#10 counter$count = 81445;
	#10 counter$count = 81446;
	#10 counter$count = 81447;
	#10 counter$count = 81448;
	#10 counter$count = 81449;
	#10 counter$count = 81450;
	#10 counter$count = 81451;
	#10 counter$count = 81452;
	#10 counter$count = 81453;
	#10 counter$count = 81454;
	#10 counter$count = 81455;
	#10 counter$count = 81456;
	#10 counter$count = 81457;
	#10 counter$count = 81458;
	#10 counter$count = 81459;
	#10 counter$count = 81460;
	#10 counter$count = 81461;
	#10 counter$count = 81462;
	#10 counter$count = 81463;
	#10 counter$count = 81464;
	#10 counter$count = 81465;
	#10 counter$count = 81466;
	#10 counter$count = 81467;
	#10 counter$count = 81468;
	#10 counter$count = 81469;
	#10 counter$count = 81470;
	#10 counter$count = 81471;
	#10 counter$count = 81472;
	#10 counter$count = 81473;
	#10 counter$count = 81474;
	#10 counter$count = 81475;
	#10 counter$count = 81476;
	#10 counter$count = 81477;
	#10 counter$count = 81478;
	#10 counter$count = 81479;
	#10 counter$count = 81480;
	#10 counter$count = 81481;
	#10 counter$count = 81482;
	#10 counter$count = 81483;
	#10 counter$count = 81484;
	#10 counter$count = 81485;
	#10 counter$count = 81486;
	#10 counter$count = 81487;
	#10 counter$count = 81488;
	#10 counter$count = 81489;
	#10 counter$count = 81490;
	#10 counter$count = 81491;
	#10 counter$count = 81492;
	#10 counter$count = 81493;
	#10 counter$count = 81494;
	#10 counter$count = 81495;
	#10 counter$count = 81496;
	#10 counter$count = 81497;
	#10 counter$count = 81498;
	#10 counter$count = 81499;
	#10 counter$count = 81500;
	#10 counter$count = 81501;
	#10 counter$count = 81502;
	#10 counter$count = 81503;
	#10 counter$count = 81504;
	#10 counter$count = 81505;
	#10 counter$count = 81506;
	#10 counter$count = 81507;
	#10 counter$count = 81508;
	#10 counter$count = 81509;
	#10 counter$count = 81510;
	#10 counter$count = 81511;
	#10 counter$count = 81512;
	#10 counter$count = 81513;
	#10 counter$count = 81514;
	#10 counter$count = 81515;
	#10 counter$count = 81516;
	#10 counter$count = 81517;
	#10 counter$count = 81518;
	#10 counter$count = 81519;
	#10 counter$count = 81520;
	#10 counter$count = 81521;
	#10 counter$count = 81522;
	#10 counter$count = 81523;
	#10 counter$count = 81524;
	#10 counter$count = 81525;
	#10 counter$count = 81526;
	#10 counter$count = 81527;
	#10 counter$count = 81528;
	#10 counter$count = 81529;
	#10 counter$count = 81530;
	#10 counter$count = 81531;
	#10 counter$count = 81532;
	#10 counter$count = 81533;
	#10 counter$count = 81534;
	#10 counter$count = 81535;
	#10 counter$count = 81536;
	#10 counter$count = 81537;
	#10 counter$count = 81538;
	#10 counter$count = 81539;
	#10 counter$count = 81540;
	#10 counter$count = 81541;
	#10 counter$count = 81542;
	#10 counter$count = 81543;
	#10 counter$count = 81544;
	#10 counter$count = 81545;
	#10 counter$count = 81546;
	#10 counter$count = 81547;
	#10 counter$count = 81548;
	#10 counter$count = 81549;
	#10 counter$count = 81550;
	#10 counter$count = 81551;
	#10 counter$count = 81552;
	#10 counter$count = 81553;
	#10 counter$count = 81554;
	#10 counter$count = 81555;
	#10 counter$count = 81556;
	#10 counter$count = 81557;
	#10 counter$count = 81558;
	#10 counter$count = 81559;
	#10 counter$count = 81560;
	#10 counter$count = 81561;
	#10 counter$count = 81562;
	#10 counter$count = 81563;
	#10 counter$count = 81564;
	#10 counter$count = 81565;
	#10 counter$count = 81566;
	#10 counter$count = 81567;
	#10 counter$count = 81568;
	#10 counter$count = 81569;
	#10 counter$count = 81570;
	#10 counter$count = 81571;
	#10 counter$count = 81572;
	#10 counter$count = 81573;
	#10 counter$count = 81574;
	#10 counter$count = 81575;
	#10 counter$count = 81576;
	#10 counter$count = 81577;
	#10 counter$count = 81578;
	#10 counter$count = 81579;
	#10 counter$count = 81580;
	#10 counter$count = 81581;
	#10 counter$count = 81582;
	#10 counter$count = 81583;
	#10 counter$count = 81584;
	#10 counter$count = 81585;
	#10 counter$count = 81586;
	#10 counter$count = 81587;
	#10 counter$count = 81588;
	#10 counter$count = 81589;
	#10 counter$count = 81590;
	#10 counter$count = 81591;
	#10 counter$count = 81592;
	#10 counter$count = 81593;
	#10 counter$count = 81594;
	#10 counter$count = 81595;
	#10 counter$count = 81596;
	#10 counter$count = 81597;
	#10 counter$count = 81598;
	#10 counter$count = 81599;
	#10 counter$count = 81600;
	#10 counter$count = 81601;
	#10 counter$count = 81602;
	#10 counter$count = 81603;
	#10 counter$count = 81604;
	#10 counter$count = 81605;
	#10 counter$count = 81606;
	#10 counter$count = 81607;
	#10 counter$count = 81608;
	#10 counter$count = 81609;
	#10 counter$count = 81610;
	#10 counter$count = 81611;
	#10 counter$count = 81612;
	#10 counter$count = 81613;
	#10 counter$count = 81614;
	#10 counter$count = 81615;
	#10 counter$count = 81616;
	#10 counter$count = 81617;
	#10 counter$count = 81618;
	#10 counter$count = 81619;
	#10 counter$count = 81620;
	#10 counter$count = 81621;
	#10 counter$count = 81622;
	#10 counter$count = 81623;
	#10 counter$count = 81624;
	#10 counter$count = 81625;
	#10 counter$count = 81626;
	#10 counter$count = 81627;
	#10 counter$count = 81628;
	#10 counter$count = 81629;
	#10 counter$count = 81630;
	#10 counter$count = 81631;
	#10 counter$count = 81632;
	#10 counter$count = 81633;
	#10 counter$count = 81634;
	#10 counter$count = 81635;
	#10 counter$count = 81636;
	#10 counter$count = 81637;
	#10 counter$count = 81638;
	#10 counter$count = 81639;
	#10 counter$count = 81640;
	#10 counter$count = 81641;
	#10 counter$count = 81642;
	#10 counter$count = 81643;
	#10 counter$count = 81644;
	#10 counter$count = 81645;
	#10 counter$count = 81646;
	#10 counter$count = 81647;
	#10 counter$count = 81648;
	#10 counter$count = 81649;
	#10 counter$count = 81650;
	#10 counter$count = 81651;
	#10 counter$count = 81652;
	#10 counter$count = 81653;
	#10 counter$count = 81654;
	#10 counter$count = 81655;
	#10 counter$count = 81656;
	#10 counter$count = 81657;
	#10 counter$count = 81658;
	#10 counter$count = 81659;
	#10 counter$count = 81660;
	#10 counter$count = 81661;
	#10 counter$count = 81662;
	#10 counter$count = 81663;
	#10 counter$count = 81664;
	#10 counter$count = 81665;
	#10 counter$count = 81666;
	#10 counter$count = 81667;
	#10 counter$count = 81668;
	#10 counter$count = 81669;
	#10 counter$count = 81670;
	#10 counter$count = 81671;
	#10 counter$count = 81672;
	#10 counter$count = 81673;
	#10 counter$count = 81674;
	#10 counter$count = 81675;
	#10 counter$count = 81676;
	#10 counter$count = 81677;
	#10 counter$count = 81678;
	#10 counter$count = 81679;
	#10 counter$count = 81680;
	#10 counter$count = 81681;
	#10 counter$count = 81682;
	#10 counter$count = 81683;
	#10 counter$count = 81684;
	#10 counter$count = 81685;
	#10 counter$count = 81686;
	#10 counter$count = 81687;
	#10 counter$count = 81688;
	#10 counter$count = 81689;
	#10 counter$count = 81690;
	#10 counter$count = 81691;
	#10 counter$count = 81692;
	#10 counter$count = 81693;
	#10 counter$count = 81694;
	#10 counter$count = 81695;
	#10 counter$count = 81696;
	#10 counter$count = 81697;
	#10 counter$count = 81698;
	#10 counter$count = 81699;
	#10 counter$count = 81700;
	#10 counter$count = 81701;
	#10 counter$count = 81702;
	#10 counter$count = 81703;
	#10 counter$count = 81704;
	#10 counter$count = 81705;
	#10 counter$count = 81706;
	#10 counter$count = 81707;
	#10 counter$count = 81708;
	#10 counter$count = 81709;
	#10 counter$count = 81710;
	#10 counter$count = 81711;
	#10 counter$count = 81712;
	#10 counter$count = 81713;
	#10 counter$count = 81714;
	#10 counter$count = 81715;
	#10 counter$count = 81716;
	#10 counter$count = 81717;
	#10 counter$count = 81718;
	#10 counter$count = 81719;
	#10 counter$count = 81720;
	#10 counter$count = 81721;
	#10 counter$count = 81722;
	#10 counter$count = 81723;
	#10 counter$count = 81724;
	#10 counter$count = 81725;
	#10 counter$count = 81726;
	#10 counter$count = 81727;
	#10 counter$count = 81728;
	#10 counter$count = 81729;
	#10 counter$count = 81730;
	#10 counter$count = 81731;
	#10 counter$count = 81732;
	#10 counter$count = 81733;
	#10 counter$count = 81734;
	#10 counter$count = 81735;
	#10 counter$count = 81736;
	#10 counter$count = 81737;
	#10 counter$count = 81738;
	#10 counter$count = 81739;
	#10 counter$count = 81740;
	#10 counter$count = 81741;
	#10 counter$count = 81742;
	#10 counter$count = 81743;
	#10 counter$count = 81744;
	#10 counter$count = 81745;
	#10 counter$count = 81746;
	#10 counter$count = 81747;
	#10 counter$count = 81748;
	#10 counter$count = 81749;
	#10 counter$count = 81750;
	#10 counter$count = 81751;
	#10 counter$count = 81752;
	#10 counter$count = 81753;
	#10 counter$count = 81754;
	#10 counter$count = 81755;
	#10 counter$count = 81756;
	#10 counter$count = 81757;
	#10 counter$count = 81758;
	#10 counter$count = 81759;
	#10 counter$count = 81760;
	#10 counter$count = 81761;
	#10 counter$count = 81762;
	#10 counter$count = 81763;
	#10 counter$count = 81764;
	#10 counter$count = 81765;
	#10 counter$count = 81766;
	#10 counter$count = 81767;
	#10 counter$count = 81768;
	#10 counter$count = 81769;
	#10 counter$count = 81770;
	#10 counter$count = 81771;
	#10 counter$count = 81772;
	#10 counter$count = 81773;
	#10 counter$count = 81774;
	#10 counter$count = 81775;
	#10 counter$count = 81776;
	#10 counter$count = 81777;
	#10 counter$count = 81778;
	#10 counter$count = 81779;
	#10 counter$count = 81780;
	#10 counter$count = 81781;
	#10 counter$count = 81782;
	#10 counter$count = 81783;
	#10 counter$count = 81784;
	#10 counter$count = 81785;
	#10 counter$count = 81786;
	#10 counter$count = 81787;
	#10 counter$count = 81788;
	#10 counter$count = 81789;
	#10 counter$count = 81790;
	#10 counter$count = 81791;
	#10 counter$count = 81792;
	#10 counter$count = 81793;
	#10 counter$count = 81794;
	#10 counter$count = 81795;
	#10 counter$count = 81796;
	#10 counter$count = 81797;
	#10 counter$count = 81798;
	#10 counter$count = 81799;
	#10 counter$count = 81800;
	#10 counter$count = 81801;
	#10 counter$count = 81802;
	#10 counter$count = 81803;
	#10 counter$count = 81804;
	#10 counter$count = 81805;
	#10 counter$count = 81806;
	#10 counter$count = 81807;
	#10 counter$count = 81808;
	#10 counter$count = 81809;
	#10 counter$count = 81810;
	#10 counter$count = 81811;
	#10 counter$count = 81812;
	#10 counter$count = 81813;
	#10 counter$count = 81814;
	#10 counter$count = 81815;
	#10 counter$count = 81816;
	#10 counter$count = 81817;
	#10 counter$count = 81818;
	#10 counter$count = 81819;
	#10 counter$count = 81820;
	#10 counter$count = 81821;
	#10 counter$count = 81822;
	#10 counter$count = 81823;
	#10 counter$count = 81824;
	#10 counter$count = 81825;
	#10 counter$count = 81826;
	#10 counter$count = 81827;
	#10 counter$count = 81828;
	#10 counter$count = 81829;
	#10 counter$count = 81830;
	#10 counter$count = 81831;
	#10 counter$count = 81832;
	#10 counter$count = 81833;
	#10 counter$count = 81834;
	#10 counter$count = 81835;
	#10 counter$count = 81836;
	#10 counter$count = 81837;
	#10 counter$count = 81838;
	#10 counter$count = 81839;
	#10 counter$count = 81840;
	#10 counter$count = 81841;
	#10 counter$count = 81842;
	#10 counter$count = 81843;
	#10 counter$count = 81844;
	#10 counter$count = 81845;
	#10 counter$count = 81846;
	#10 counter$count = 81847;
	#10 counter$count = 81848;
	#10 counter$count = 81849;
	#10 counter$count = 81850;
	#10 counter$count = 81851;
	#10 counter$count = 81852;
	#10 counter$count = 81853;
	#10 counter$count = 81854;
	#10 counter$count = 81855;
	#10 counter$count = 81856;
	#10 counter$count = 81857;
	#10 counter$count = 81858;
	#10 counter$count = 81859;
	#10 counter$count = 81860;
	#10 counter$count = 81861;
	#10 counter$count = 81862;
	#10 counter$count = 81863;
	#10 counter$count = 81864;
	#10 counter$count = 81865;
	#10 counter$count = 81866;
	#10 counter$count = 81867;
	#10 counter$count = 81868;
	#10 counter$count = 81869;
	#10 counter$count = 81870;
	#10 counter$count = 81871;
	#10 counter$count = 81872;
	#10 counter$count = 81873;
	#10 counter$count = 81874;
	#10 counter$count = 81875;
	#10 counter$count = 81876;
	#10 counter$count = 81877;
	#10 counter$count = 81878;
	#10 counter$count = 81879;
	#10 counter$count = 81880;
	#10 counter$count = 81881;
	#10 counter$count = 81882;
	#10 counter$count = 81883;
	#10 counter$count = 81884;
	#10 counter$count = 81885;
	#10 counter$count = 81886;
	#10 counter$count = 81887;
	#10 counter$count = 81888;
	#10 counter$count = 81889;
	#10 counter$count = 81890;
	#10 counter$count = 81891;
	#10 counter$count = 81892;
	#10 counter$count = 81893;
	#10 counter$count = 81894;
	#10 counter$count = 81895;
	#10 counter$count = 81896;
	#10 counter$count = 81897;
	#10 counter$count = 81898;
	#10 counter$count = 81899;
	#10 counter$count = 81900;
	#10 counter$count = 81901;
	#10 counter$count = 81902;
	#10 counter$count = 81903;
	#10 counter$count = 81904;
	#10 counter$count = 81905;
	#10 counter$count = 81906;
	#10 counter$count = 81907;
	#10 counter$count = 81908;
	#10 counter$count = 81909;
	#10 counter$count = 81910;
	#10 counter$count = 81911;
	#10 counter$count = 81912;
	#10 counter$count = 81913;
	#10 counter$count = 81914;
	#10 counter$count = 81915;
	#10 counter$count = 81916;
	#10 counter$count = 81917;
	#10 counter$count = 81918;
	#10 counter$count = 81919;
	#10 counter$count = 81920;
	#10 counter$count = 81921;
	#10 counter$count = 81922;
	#10 counter$count = 81923;
	#10 counter$count = 81924;
	#10 counter$count = 81925;
	#10 counter$count = 81926;
	#10 counter$count = 81927;
	#10 counter$count = 81928;
	#10 counter$count = 81929;
	#10 counter$count = 81930;
	#10 counter$count = 81931;
	#10 counter$count = 81932;
	#10 counter$count = 81933;
	#10 counter$count = 81934;
	#10 counter$count = 81935;
	#10 counter$count = 81936;
	#10 counter$count = 81937;
	#10 counter$count = 81938;
	#10 counter$count = 81939;
	#10 counter$count = 81940;
	#10 counter$count = 81941;
	#10 counter$count = 81942;
	#10 counter$count = 81943;
	#10 counter$count = 81944;
	#10 counter$count = 81945;
	#10 counter$count = 81946;
	#10 counter$count = 81947;
	#10 counter$count = 81948;
	#10 counter$count = 81949;
	#10 counter$count = 81950;
	#10 counter$count = 81951;
	#10 counter$count = 81952;
	#10 counter$count = 81953;
	#10 counter$count = 81954;
	#10 counter$count = 81955;
	#10 counter$count = 81956;
	#10 counter$count = 81957;
	#10 counter$count = 81958;
	#10 counter$count = 81959;
	#10 counter$count = 81960;
	#10 counter$count = 81961;
	#10 counter$count = 81962;
	#10 counter$count = 81963;
	#10 counter$count = 81964;
	#10 counter$count = 81965;
	#10 counter$count = 81966;
	#10 counter$count = 81967;
	#10 counter$count = 81968;
	#10 counter$count = 81969;
	#10 counter$count = 81970;
	#10 counter$count = 81971;
	#10 counter$count = 81972;
	#10 counter$count = 81973;
	#10 counter$count = 81974;
	#10 counter$count = 81975;
	#10 counter$count = 81976;
	#10 counter$count = 81977;
	#10 counter$count = 81978;
	#10 counter$count = 81979;
	#10 counter$count = 81980;
	#10 counter$count = 81981;
	#10 counter$count = 81982;
	#10 counter$count = 81983;
	#10 counter$count = 81984;
	#10 counter$count = 81985;
	#10 counter$count = 81986;
	#10 counter$count = 81987;
	#10 counter$count = 81988;
	#10 counter$count = 81989;
	#10 counter$count = 81990;
	#10 counter$count = 81991;
	#10 counter$count = 81992;
	#10 counter$count = 81993;
	#10 counter$count = 81994;
	#10 counter$count = 81995;
	#10 counter$count = 81996;
	#10 counter$count = 81997;
	#10 counter$count = 81998;
	#10 counter$count = 81999;
	#10 counter$count = 82000;
	#10 counter$count = 82001;
	#10 counter$count = 82002;
	#10 counter$count = 82003;
	#10 counter$count = 82004;
	#10 counter$count = 82005;
	#10 counter$count = 82006;
	#10 counter$count = 82007;
	#10 counter$count = 82008;
	#10 counter$count = 82009;
	#10 counter$count = 82010;
	#10 counter$count = 82011;
	#10 counter$count = 82012;
	#10 counter$count = 82013;
	#10 counter$count = 82014;
	#10 counter$count = 82015;
	#10 counter$count = 82016;
	#10 counter$count = 82017;
	#10 counter$count = 82018;
	#10 counter$count = 82019;
	#10 counter$count = 82020;
	#10 counter$count = 82021;
	#10 counter$count = 82022;
	#10 counter$count = 82023;
	#10 counter$count = 82024;
	#10 counter$count = 82025;
	#10 counter$count = 82026;
	#10 counter$count = 82027;
	#10 counter$count = 82028;
	#10 counter$count = 82029;
	#10 counter$count = 82030;
	#10 counter$count = 82031;
	#10 counter$count = 82032;
	#10 counter$count = 82033;
	#10 counter$count = 82034;
	#10 counter$count = 82035;
	#10 counter$count = 82036;
	#10 counter$count = 82037;
	#10 counter$count = 82038;
	#10 counter$count = 82039;
	#10 counter$count = 82040;
	#10 counter$count = 82041;
	#10 counter$count = 82042;
	#10 counter$count = 82043;
	#10 counter$count = 82044;
	#10 counter$count = 82045;
	#10 counter$count = 82046;
	#10 counter$count = 82047;
	#10 counter$count = 82048;
	#10 counter$count = 82049;
	#10 counter$count = 82050;
	#10 counter$count = 82051;
	#10 counter$count = 82052;
	#10 counter$count = 82053;
	#10 counter$count = 82054;
	#10 counter$count = 82055;
	#10 counter$count = 82056;
	#10 counter$count = 82057;
	#10 counter$count = 82058;
	#10 counter$count = 82059;
	#10 counter$count = 82060;
	#10 counter$count = 82061;
	#10 counter$count = 82062;
	#10 counter$count = 82063;
	#10 counter$count = 82064;
	#10 counter$count = 82065;
	#10 counter$count = 82066;
	#10 counter$count = 82067;
	#10 counter$count = 82068;
	#10 counter$count = 82069;
	#10 counter$count = 82070;
	#10 counter$count = 82071;
	#10 counter$count = 82072;
	#10 counter$count = 82073;
	#10 counter$count = 82074;
	#10 counter$count = 82075;
	#10 counter$count = 82076;
	#10 counter$count = 82077;
	#10 counter$count = 82078;
	#10 counter$count = 82079;
	#10 counter$count = 82080;
	#10 counter$count = 82081;
	#10 counter$count = 82082;
	#10 counter$count = 82083;
	#10 counter$count = 82084;
	#10 counter$count = 82085;
	#10 counter$count = 82086;
	#10 counter$count = 82087;
	#10 counter$count = 82088;
	#10 counter$count = 82089;
	#10 counter$count = 82090;
	#10 counter$count = 82091;
	#10 counter$count = 82092;
	#10 counter$count = 82093;
	#10 counter$count = 82094;
	#10 counter$count = 82095;
	#10 counter$count = 82096;
	#10 counter$count = 82097;
	#10 counter$count = 82098;
	#10 counter$count = 82099;
	#10 counter$count = 82100;
	#10 counter$count = 82101;
	#10 counter$count = 82102;
	#10 counter$count = 82103;
	#10 counter$count = 82104;
	#10 counter$count = 82105;
	#10 counter$count = 82106;
	#10 counter$count = 82107;
	#10 counter$count = 82108;
	#10 counter$count = 82109;
	#10 counter$count = 82110;
	#10 counter$count = 82111;
	#10 counter$count = 82112;
	#10 counter$count = 82113;
	#10 counter$count = 82114;
	#10 counter$count = 82115;
	#10 counter$count = 82116;
	#10 counter$count = 82117;
	#10 counter$count = 82118;
	#10 counter$count = 82119;
	#10 counter$count = 82120;
	#10 counter$count = 82121;
	#10 counter$count = 82122;
	#10 counter$count = 82123;
	#10 counter$count = 82124;
	#10 counter$count = 82125;
	#10 counter$count = 82126;
	#10 counter$count = 82127;
	#10 counter$count = 82128;
	#10 counter$count = 82129;
	#10 counter$count = 82130;
	#10 counter$count = 82131;
	#10 counter$count = 82132;
	#10 counter$count = 82133;
	#10 counter$count = 82134;
	#10 counter$count = 82135;
	#10 counter$count = 82136;
	#10 counter$count = 82137;
	#10 counter$count = 82138;
	#10 counter$count = 82139;
	#10 counter$count = 82140;
	#10 counter$count = 82141;
	#10 counter$count = 82142;
	#10 counter$count = 82143;
	#10 counter$count = 82144;
	#10 counter$count = 82145;
	#10 counter$count = 82146;
	#10 counter$count = 82147;
	#10 counter$count = 82148;
	#10 counter$count = 82149;
	#10 counter$count = 82150;
	#10 counter$count = 82151;
	#10 counter$count = 82152;
	#10 counter$count = 82153;
	#10 counter$count = 82154;
	#10 counter$count = 82155;
	#10 counter$count = 82156;
	#10 counter$count = 82157;
	#10 counter$count = 82158;
	#10 counter$count = 82159;
	#10 counter$count = 82160;
	#10 counter$count = 82161;
	#10 counter$count = 82162;
	#10 counter$count = 82163;
	#10 counter$count = 82164;
	#10 counter$count = 82165;
	#10 counter$count = 82166;
	#10 counter$count = 82167;
	#10 counter$count = 82168;
	#10 counter$count = 82169;
	#10 counter$count = 82170;
	#10 counter$count = 82171;
	#10 counter$count = 82172;
	#10 counter$count = 82173;
	#10 counter$count = 82174;
	#10 counter$count = 82175;
	#10 counter$count = 82176;
	#10 counter$count = 82177;
	#10 counter$count = 82178;
	#10 counter$count = 82179;
	#10 counter$count = 82180;
	#10 counter$count = 82181;
	#10 counter$count = 82182;
	#10 counter$count = 82183;
	#10 counter$count = 82184;
	#10 counter$count = 82185;
	#10 counter$count = 82186;
	#10 counter$count = 82187;
	#10 counter$count = 82188;
	#10 counter$count = 82189;
	#10 counter$count = 82190;
	#10 counter$count = 82191;
	#10 counter$count = 82192;
	#10 counter$count = 82193;
	#10 counter$count = 82194;
	#10 counter$count = 82195;
	#10 counter$count = 82196;
	#10 counter$count = 82197;
	#10 counter$count = 82198;
	#10 counter$count = 82199;
	#10 counter$count = 82200;
	#10 counter$count = 82201;
	#10 counter$count = 82202;
	#10 counter$count = 82203;
	#10 counter$count = 82204;
	#10 counter$count = 82205;
	#10 counter$count = 82206;
	#10 counter$count = 82207;
	#10 counter$count = 82208;
	#10 counter$count = 82209;
	#10 counter$count = 82210;
	#10 counter$count = 82211;
	#10 counter$count = 82212;
	#10 counter$count = 82213;
	#10 counter$count = 82214;
	#10 counter$count = 82215;
	#10 counter$count = 82216;
	#10 counter$count = 82217;
	#10 counter$count = 82218;
	#10 counter$count = 82219;
	#10 counter$count = 82220;
	#10 counter$count = 82221;
	#10 counter$count = 82222;
	#10 counter$count = 82223;
	#10 counter$count = 82224;
	#10 counter$count = 82225;
	#10 counter$count = 82226;
	#10 counter$count = 82227;
	#10 counter$count = 82228;
	#10 counter$count = 82229;
	#10 counter$count = 82230;
	#10 counter$count = 82231;
	#10 counter$count = 82232;
	#10 counter$count = 82233;
	#10 counter$count = 82234;
	#10 counter$count = 82235;
	#10 counter$count = 82236;
	#10 counter$count = 82237;
	#10 counter$count = 82238;
	#10 counter$count = 82239;
	#10 counter$count = 82240;
	#10 counter$count = 82241;
	#10 counter$count = 82242;
	#10 counter$count = 82243;
	#10 counter$count = 82244;
	#10 counter$count = 82245;
	#10 counter$count = 82246;
	#10 counter$count = 82247;
	#10 counter$count = 82248;
	#10 counter$count = 82249;
	#10 counter$count = 82250;
	#10 counter$count = 82251;
	#10 counter$count = 82252;
	#10 counter$count = 82253;
	#10 counter$count = 82254;
	#10 counter$count = 82255;
	#10 counter$count = 82256;
	#10 counter$count = 82257;
	#10 counter$count = 82258;
	#10 counter$count = 82259;
	#10 counter$count = 82260;
	#10 counter$count = 82261;
	#10 counter$count = 82262;
	#10 counter$count = 82263;
	#10 counter$count = 82264;
	#10 counter$count = 82265;
	#10 counter$count = 82266;
	#10 counter$count = 82267;
	#10 counter$count = 82268;
	#10 counter$count = 82269;
	#10 counter$count = 82270;
	#10 counter$count = 82271;
	#10 counter$count = 82272;
	#10 counter$count = 82273;
	#10 counter$count = 82274;
	#10 counter$count = 82275;
	#10 counter$count = 82276;
	#10 counter$count = 82277;
	#10 counter$count = 82278;
	#10 counter$count = 82279;
	#10 counter$count = 82280;
	#10 counter$count = 82281;
	#10 counter$count = 82282;
	#10 counter$count = 82283;
	#10 counter$count = 82284;
	#10 counter$count = 82285;
	#10 counter$count = 82286;
	#10 counter$count = 82287;
	#10 counter$count = 82288;
	#10 counter$count = 82289;
	#10 counter$count = 82290;
	#10 counter$count = 82291;
	#10 counter$count = 82292;
	#10 counter$count = 82293;
	#10 counter$count = 82294;
	#10 counter$count = 82295;
	#10 counter$count = 82296;
	#10 counter$count = 82297;
	#10 counter$count = 82298;
	#10 counter$count = 82299;
	#10 counter$count = 82300;
	#10 counter$count = 82301;
	#10 counter$count = 82302;
	#10 counter$count = 82303;
	#10 counter$count = 82304;
	#10 counter$count = 82305;
	#10 counter$count = 82306;
	#10 counter$count = 82307;
	#10 counter$count = 82308;
	#10 counter$count = 82309;
	#10 counter$count = 82310;
	#10 counter$count = 82311;
	#10 counter$count = 82312;
	#10 counter$count = 82313;
	#10 counter$count = 82314;
	#10 counter$count = 82315;
	#10 counter$count = 82316;
	#10 counter$count = 82317;
	#10 counter$count = 82318;
	#10 counter$count = 82319;
	#10 counter$count = 82320;
	#10 counter$count = 82321;
	#10 counter$count = 82322;
	#10 counter$count = 82323;
	#10 counter$count = 82324;
	#10 counter$count = 82325;
	#10 counter$count = 82326;
	#10 counter$count = 82327;
	#10 counter$count = 82328;
	#10 counter$count = 82329;
	#10 counter$count = 82330;
	#10 counter$count = 82331;
	#10 counter$count = 82332;
	#10 counter$count = 82333;
	#10 counter$count = 82334;
	#10 counter$count = 82335;
	#10 counter$count = 82336;
	#10 counter$count = 82337;
	#10 counter$count = 82338;
	#10 counter$count = 82339;
	#10 counter$count = 82340;
	#10 counter$count = 82341;
	#10 counter$count = 82342;
	#10 counter$count = 82343;
	#10 counter$count = 82344;
	#10 counter$count = 82345;
	#10 counter$count = 82346;
	#10 counter$count = 82347;
	#10 counter$count = 82348;
	#10 counter$count = 82349;
	#10 counter$count = 82350;
	#10 counter$count = 82351;
	#10 counter$count = 82352;
	#10 counter$count = 82353;
	#10 counter$count = 82354;
	#10 counter$count = 82355;
	#10 counter$count = 82356;
	#10 counter$count = 82357;
	#10 counter$count = 82358;
	#10 counter$count = 82359;
	#10 counter$count = 82360;
	#10 counter$count = 82361;
	#10 counter$count = 82362;
	#10 counter$count = 82363;
	#10 counter$count = 82364;
	#10 counter$count = 82365;
	#10 counter$count = 82366;
	#10 counter$count = 82367;
	#10 counter$count = 82368;
	#10 counter$count = 82369;
	#10 counter$count = 82370;
	#10 counter$count = 82371;
	#10 counter$count = 82372;
	#10 counter$count = 82373;
	#10 counter$count = 82374;
	#10 counter$count = 82375;
	#10 counter$count = 82376;
	#10 counter$count = 82377;
	#10 counter$count = 82378;
	#10 counter$count = 82379;
	#10 counter$count = 82380;
	#10 counter$count = 82381;
	#10 counter$count = 82382;
	#10 counter$count = 82383;
	#10 counter$count = 82384;
	#10 counter$count = 82385;
	#10 counter$count = 82386;
	#10 counter$count = 82387;
	#10 counter$count = 82388;
	#10 counter$count = 82389;
	#10 counter$count = 82390;
	#10 counter$count = 82391;
	#10 counter$count = 82392;
	#10 counter$count = 82393;
	#10 counter$count = 82394;
	#10 counter$count = 82395;
	#10 counter$count = 82396;
	#10 counter$count = 82397;
	#10 counter$count = 82398;
	#10 counter$count = 82399;
	#10 counter$count = 82400;
	#10 counter$count = 82401;
	#10 counter$count = 82402;
	#10 counter$count = 82403;
	#10 counter$count = 82404;
	#10 counter$count = 82405;
	#10 counter$count = 82406;
	#10 counter$count = 82407;
	#10 counter$count = 82408;
	#10 counter$count = 82409;
	#10 counter$count = 82410;
	#10 counter$count = 82411;
	#10 counter$count = 82412;
	#10 counter$count = 82413;
	#10 counter$count = 82414;
	#10 counter$count = 82415;
	#10 counter$count = 82416;
	#10 counter$count = 82417;
	#10 counter$count = 82418;
	#10 counter$count = 82419;
	#10 counter$count = 82420;
	#10 counter$count = 82421;
	#10 counter$count = 82422;
	#10 counter$count = 82423;
	#10 counter$count = 82424;
	#10 counter$count = 82425;
	#10 counter$count = 82426;
	#10 counter$count = 82427;
	#10 counter$count = 82428;
	#10 counter$count = 82429;
	#10 counter$count = 82430;
	#10 counter$count = 82431;
	#10 counter$count = 82432;
	#10 counter$count = 82433;
	#10 counter$count = 82434;
	#10 counter$count = 82435;
	#10 counter$count = 82436;
	#10 counter$count = 82437;
	#10 counter$count = 82438;
	#10 counter$count = 82439;
	#10 counter$count = 82440;
	#10 counter$count = 82441;
	#10 counter$count = 82442;
	#10 counter$count = 82443;
	#10 counter$count = 82444;
	#10 counter$count = 82445;
	#10 counter$count = 82446;
	#10 counter$count = 82447;
	#10 counter$count = 82448;
	#10 counter$count = 82449;
	#10 counter$count = 82450;
	#10 counter$count = 82451;
	#10 counter$count = 82452;
	#10 counter$count = 82453;
	#10 counter$count = 82454;
	#10 counter$count = 82455;
	#10 counter$count = 82456;
	#10 counter$count = 82457;
	#10 counter$count = 82458;
	#10 counter$count = 82459;
	#10 counter$count = 82460;
	#10 counter$count = 82461;
	#10 counter$count = 82462;
	#10 counter$count = 82463;
	#10 counter$count = 82464;
	#10 counter$count = 82465;
	#10 counter$count = 82466;
	#10 counter$count = 82467;
	#10 counter$count = 82468;
	#10 counter$count = 82469;
	#10 counter$count = 82470;
	#10 counter$count = 82471;
	#10 counter$count = 82472;
	#10 counter$count = 82473;
	#10 counter$count = 82474;
	#10 counter$count = 82475;
	#10 counter$count = 82476;
	#10 counter$count = 82477;
	#10 counter$count = 82478;
	#10 counter$count = 82479;
	#10 counter$count = 82480;
	#10 counter$count = 82481;
	#10 counter$count = 82482;
	#10 counter$count = 82483;
	#10 counter$count = 82484;
	#10 counter$count = 82485;
	#10 counter$count = 82486;
	#10 counter$count = 82487;
	#10 counter$count = 82488;
	#10 counter$count = 82489;
	#10 counter$count = 82490;
	#10 counter$count = 82491;
	#10 counter$count = 82492;
	#10 counter$count = 82493;
	#10 counter$count = 82494;
	#10 counter$count = 82495;
	#10 counter$count = 82496;
	#10 counter$count = 82497;
	#10 counter$count = 82498;
	#10 counter$count = 82499;
	#10 counter$count = 82500;
	#10 counter$count = 82501;
	#10 counter$count = 82502;
	#10 counter$count = 82503;
	#10 counter$count = 82504;
	#10 counter$count = 82505;
	#10 counter$count = 82506;
	#10 counter$count = 82507;
	#10 counter$count = 82508;
	#10 counter$count = 82509;
	#10 counter$count = 82510;
	#10 counter$count = 82511;
	#10 counter$count = 82512;
	#10 counter$count = 82513;
	#10 counter$count = 82514;
	#10 counter$count = 82515;
	#10 counter$count = 82516;
	#10 counter$count = 82517;
	#10 counter$count = 82518;
	#10 counter$count = 82519;
	#10 counter$count = 82520;
	#10 counter$count = 82521;
	#10 counter$count = 82522;
	#10 counter$count = 82523;
	#10 counter$count = 82524;
	#10 counter$count = 82525;
	#10 counter$count = 82526;
	#10 counter$count = 82527;
	#10 counter$count = 82528;
	#10 counter$count = 82529;
	#10 counter$count = 82530;
	#10 counter$count = 82531;
	#10 counter$count = 82532;
	#10 counter$count = 82533;
	#10 counter$count = 82534;
	#10 counter$count = 82535;
	#10 counter$count = 82536;
	#10 counter$count = 82537;
	#10 counter$count = 82538;
	#10 counter$count = 82539;
	#10 counter$count = 82540;
	#10 counter$count = 82541;
	#10 counter$count = 82542;
	#10 counter$count = 82543;
	#10 counter$count = 82544;
	#10 counter$count = 82545;
	#10 counter$count = 82546;
	#10 counter$count = 82547;
	#10 counter$count = 82548;
	#10 counter$count = 82549;
	#10 counter$count = 82550;
	#10 counter$count = 82551;
	#10 counter$count = 82552;
	#10 counter$count = 82553;
	#10 counter$count = 82554;
	#10 counter$count = 82555;
	#10 counter$count = 82556;
	#10 counter$count = 82557;
	#10 counter$count = 82558;
	#10 counter$count = 82559;
	#10 counter$count = 82560;
	#10 counter$count = 82561;
	#10 counter$count = 82562;
	#10 counter$count = 82563;
	#10 counter$count = 82564;
	#10 counter$count = 82565;
	#10 counter$count = 82566;
	#10 counter$count = 82567;
	#10 counter$count = 82568;
	#10 counter$count = 82569;
	#10 counter$count = 82570;
	#10 counter$count = 82571;
	#10 counter$count = 82572;
	#10 counter$count = 82573;
	#10 counter$count = 82574;
	#10 counter$count = 82575;
	#10 counter$count = 82576;
	#10 counter$count = 82577;
	#10 counter$count = 82578;
	#10 counter$count = 82579;
	#10 counter$count = 82580;
	#10 counter$count = 82581;
	#10 counter$count = 82582;
	#10 counter$count = 82583;
	#10 counter$count = 82584;
	#10 counter$count = 82585;
	#10 counter$count = 82586;
	#10 counter$count = 82587;
	#10 counter$count = 82588;
	#10 counter$count = 82589;
	#10 counter$count = 82590;
	#10 counter$count = 82591;
	#10 counter$count = 82592;
	#10 counter$count = 82593;
	#10 counter$count = 82594;
	#10 counter$count = 82595;
	#10 counter$count = 82596;
	#10 counter$count = 82597;
	#10 counter$count = 82598;
	#10 counter$count = 82599;
	#10 counter$count = 82600;
	#10 counter$count = 82601;
	#10 counter$count = 82602;
	#10 counter$count = 82603;
	#10 counter$count = 82604;
	#10 counter$count = 82605;
	#10 counter$count = 82606;
	#10 counter$count = 82607;
	#10 counter$count = 82608;
	#10 counter$count = 82609;
	#10 counter$count = 82610;
	#10 counter$count = 82611;
	#10 counter$count = 82612;
	#10 counter$count = 82613;
	#10 counter$count = 82614;
	#10 counter$count = 82615;
	#10 counter$count = 82616;
	#10 counter$count = 82617;
	#10 counter$count = 82618;
	#10 counter$count = 82619;
	#10 counter$count = 82620;
	#10 counter$count = 82621;
	#10 counter$count = 82622;
	#10 counter$count = 82623;
	#10 counter$count = 82624;
	#10 counter$count = 82625;
	#10 counter$count = 82626;
	#10 counter$count = 82627;
	#10 counter$count = 82628;
	#10 counter$count = 82629;
	#10 counter$count = 82630;
	#10 counter$count = 82631;
	#10 counter$count = 82632;
	#10 counter$count = 82633;
	#10 counter$count = 82634;
	#10 counter$count = 82635;
	#10 counter$count = 82636;
	#10 counter$count = 82637;
	#10 counter$count = 82638;
	#10 counter$count = 82639;
	#10 counter$count = 82640;
	#10 counter$count = 82641;
	#10 counter$count = 82642;
	#10 counter$count = 82643;
	#10 counter$count = 82644;
	#10 counter$count = 82645;
	#10 counter$count = 82646;
	#10 counter$count = 82647;
	#10 counter$count = 82648;
	#10 counter$count = 82649;
	#10 counter$count = 82650;
	#10 counter$count = 82651;
	#10 counter$count = 82652;
	#10 counter$count = 82653;
	#10 counter$count = 82654;
	#10 counter$count = 82655;
	#10 counter$count = 82656;
	#10 counter$count = 82657;
	#10 counter$count = 82658;
	#10 counter$count = 82659;
	#10 counter$count = 82660;
	#10 counter$count = 82661;
	#10 counter$count = 82662;
	#10 counter$count = 82663;
	#10 counter$count = 82664;
	#10 counter$count = 82665;
	#10 counter$count = 82666;
	#10 counter$count = 82667;
	#10 counter$count = 82668;
	#10 counter$count = 82669;
	#10 counter$count = 82670;
	#10 counter$count = 82671;
	#10 counter$count = 82672;
	#10 counter$count = 82673;
	#10 counter$count = 82674;
	#10 counter$count = 82675;
	#10 counter$count = 82676;
	#10 counter$count = 82677;
	#10 counter$count = 82678;
	#10 counter$count = 82679;
	#10 counter$count = 82680;
	#10 counter$count = 82681;
	#10 counter$count = 82682;
	#10 counter$count = 82683;
	#10 counter$count = 82684;
	#10 counter$count = 82685;
	#10 counter$count = 82686;
	#10 counter$count = 82687;
	#10 counter$count = 82688;
	#10 counter$count = 82689;
	#10 counter$count = 82690;
	#10 counter$count = 82691;
	#10 counter$count = 82692;
	#10 counter$count = 82693;
	#10 counter$count = 82694;
	#10 counter$count = 82695;
	#10 counter$count = 82696;
	#10 counter$count = 82697;
	#10 counter$count = 82698;
	#10 counter$count = 82699;
	#10 counter$count = 82700;
	#10 counter$count = 82701;
	#10 counter$count = 82702;
	#10 counter$count = 82703;
	#10 counter$count = 82704;
	#10 counter$count = 82705;
	#10 counter$count = 82706;
	#10 counter$count = 82707;
	#10 counter$count = 82708;
	#10 counter$count = 82709;
	#10 counter$count = 82710;
	#10 counter$count = 82711;
	#10 counter$count = 82712;
	#10 counter$count = 82713;
	#10 counter$count = 82714;
	#10 counter$count = 82715;
	#10 counter$count = 82716;
	#10 counter$count = 82717;
	#10 counter$count = 82718;
	#10 counter$count = 82719;
	#10 counter$count = 82720;
	#10 counter$count = 82721;
	#10 counter$count = 82722;
	#10 counter$count = 82723;
	#10 counter$count = 82724;
	#10 counter$count = 82725;
	#10 counter$count = 82726;
	#10 counter$count = 82727;
	#10 counter$count = 82728;
	#10 counter$count = 82729;
	#10 counter$count = 82730;
	#10 counter$count = 82731;
	#10 counter$count = 82732;
	#10 counter$count = 82733;
	#10 counter$count = 82734;
	#10 counter$count = 82735;
	#10 counter$count = 82736;
	#10 counter$count = 82737;
	#10 counter$count = 82738;
	#10 counter$count = 82739;
	#10 counter$count = 82740;
	#10 counter$count = 82741;
	#10 counter$count = 82742;
	#10 counter$count = 82743;
	#10 counter$count = 82744;
	#10 counter$count = 82745;
	#10 counter$count = 82746;
	#10 counter$count = 82747;
	#10 counter$count = 82748;
	#10 counter$count = 82749;
	#10 counter$count = 82750;
	#10 counter$count = 82751;
	#10 counter$count = 82752;
	#10 counter$count = 82753;
	#10 counter$count = 82754;
	#10 counter$count = 82755;
	#10 counter$count = 82756;
	#10 counter$count = 82757;
	#10 counter$count = 82758;
	#10 counter$count = 82759;
	#10 counter$count = 82760;
	#10 counter$count = 82761;
	#10 counter$count = 82762;
	#10 counter$count = 82763;
	#10 counter$count = 82764;
	#10 counter$count = 82765;
	#10 counter$count = 82766;
	#10 counter$count = 82767;
	#10 counter$count = 82768;
	#10 counter$count = 82769;
	#10 counter$count = 82770;
	#10 counter$count = 82771;
	#10 counter$count = 82772;
	#10 counter$count = 82773;
	#10 counter$count = 82774;
	#10 counter$count = 82775;
	#10 counter$count = 82776;
	#10 counter$count = 82777;
	#10 counter$count = 82778;
	#10 counter$count = 82779;
	#10 counter$count = 82780;
	#10 counter$count = 82781;
	#10 counter$count = 82782;
	#10 counter$count = 82783;
	#10 counter$count = 82784;
	#10 counter$count = 82785;
	#10 counter$count = 82786;
	#10 counter$count = 82787;
	#10 counter$count = 82788;
	#10 counter$count = 82789;
	#10 counter$count = 82790;
	#10 counter$count = 82791;
	#10 counter$count = 82792;
	#10 counter$count = 82793;
	#10 counter$count = 82794;
	#10 counter$count = 82795;
	#10 counter$count = 82796;
	#10 counter$count = 82797;
	#10 counter$count = 82798;
	#10 counter$count = 82799;
	#10 counter$count = 82800;
	#10 counter$count = 82801;
	#10 counter$count = 82802;
	#10 counter$count = 82803;
	#10 counter$count = 82804;
	#10 counter$count = 82805;
	#10 counter$count = 82806;
	#10 counter$count = 82807;
	#10 counter$count = 82808;
	#10 counter$count = 82809;
	#10 counter$count = 82810;
	#10 counter$count = 82811;
	#10 counter$count = 82812;
	#10 counter$count = 82813;
	#10 counter$count = 82814;
	#10 counter$count = 82815;
	#10 counter$count = 82816;
	#10 counter$count = 82817;
	#10 counter$count = 82818;
	#10 counter$count = 82819;
	#10 counter$count = 82820;
	#10 counter$count = 82821;
	#10 counter$count = 82822;
	#10 counter$count = 82823;
	#10 counter$count = 82824;
	#10 counter$count = 82825;
	#10 counter$count = 82826;
	#10 counter$count = 82827;
	#10 counter$count = 82828;
	#10 counter$count = 82829;
	#10 counter$count = 82830;
	#10 counter$count = 82831;
	#10 counter$count = 82832;
	#10 counter$count = 82833;
	#10 counter$count = 82834;
	#10 counter$count = 82835;
	#10 counter$count = 82836;
	#10 counter$count = 82837;
	#10 counter$count = 82838;
	#10 counter$count = 82839;
	#10 counter$count = 82840;
	#10 counter$count = 82841;
	#10 counter$count = 82842;
	#10 counter$count = 82843;
	#10 counter$count = 82844;
	#10 counter$count = 82845;
	#10 counter$count = 82846;
	#10 counter$count = 82847;
	#10 counter$count = 82848;
	#10 counter$count = 82849;
	#10 counter$count = 82850;
	#10 counter$count = 82851;
	#10 counter$count = 82852;
	#10 counter$count = 82853;
	#10 counter$count = 82854;
	#10 counter$count = 82855;
	#10 counter$count = 82856;
	#10 counter$count = 82857;
	#10 counter$count = 82858;
	#10 counter$count = 82859;
	#10 counter$count = 82860;
	#10 counter$count = 82861;
	#10 counter$count = 82862;
	#10 counter$count = 82863;
	#10 counter$count = 82864;
	#10 counter$count = 82865;
	#10 counter$count = 82866;
	#10 counter$count = 82867;
	#10 counter$count = 82868;
	#10 counter$count = 82869;
	#10 counter$count = 82870;
	#10 counter$count = 82871;
	#10 counter$count = 82872;
	#10 counter$count = 82873;
	#10 counter$count = 82874;
	#10 counter$count = 82875;
	#10 counter$count = 82876;
	#10 counter$count = 82877;
	#10 counter$count = 82878;
	#10 counter$count = 82879;
	#10 counter$count = 82880;
	#10 counter$count = 82881;
	#10 counter$count = 82882;
	#10 counter$count = 82883;
	#10 counter$count = 82884;
	#10 counter$count = 82885;
	#10 counter$count = 82886;
	#10 counter$count = 82887;
	#10 counter$count = 82888;
	#10 counter$count = 82889;
	#10 counter$count = 82890;
	#10 counter$count = 82891;
	#10 counter$count = 82892;
	#10 counter$count = 82893;
	#10 counter$count = 82894;
	#10 counter$count = 82895;
	#10 counter$count = 82896;
	#10 counter$count = 82897;
	#10 counter$count = 82898;
	#10 counter$count = 82899;
	#10 counter$count = 82900;
	#10 counter$count = 82901;
	#10 counter$count = 82902;
	#10 counter$count = 82903;
	#10 counter$count = 82904;
	#10 counter$count = 82905;
	#10 counter$count = 82906;
	#10 counter$count = 82907;
	#10 counter$count = 82908;
	#10 counter$count = 82909;
	#10 counter$count = 82910;
	#10 counter$count = 82911;
	#10 counter$count = 82912;
	#10 counter$count = 82913;
	#10 counter$count = 82914;
	#10 counter$count = 82915;
	#10 counter$count = 82916;
	#10 counter$count = 82917;
	#10 counter$count = 82918;
	#10 counter$count = 82919;
	#10 counter$count = 82920;
	#10 counter$count = 82921;
	#10 counter$count = 82922;
	#10 counter$count = 82923;
	#10 counter$count = 82924;
	#10 counter$count = 82925;
	#10 counter$count = 82926;
	#10 counter$count = 82927;
	#10 counter$count = 82928;
	#10 counter$count = 82929;
	#10 counter$count = 82930;
	#10 counter$count = 82931;
	#10 counter$count = 82932;
	#10 counter$count = 82933;
	#10 counter$count = 82934;
	#10 counter$count = 82935;
	#10 counter$count = 82936;
	#10 counter$count = 82937;
	#10 counter$count = 82938;
	#10 counter$count = 82939;
	#10 counter$count = 82940;
	#10 counter$count = 82941;
	#10 counter$count = 82942;
	#10 counter$count = 82943;
	#10 counter$count = 82944;
	#10 counter$count = 82945;
	#10 counter$count = 82946;
	#10 counter$count = 82947;
	#10 counter$count = 82948;
	#10 counter$count = 82949;
	#10 counter$count = 82950;
	#10 counter$count = 82951;
	#10 counter$count = 82952;
	#10 counter$count = 82953;
	#10 counter$count = 82954;
	#10 counter$count = 82955;
	#10 counter$count = 82956;
	#10 counter$count = 82957;
	#10 counter$count = 82958;
	#10 counter$count = 82959;
	#10 counter$count = 82960;
	#10 counter$count = 82961;
	#10 counter$count = 82962;
	#10 counter$count = 82963;
	#10 counter$count = 82964;
	#10 counter$count = 82965;
	#10 counter$count = 82966;
	#10 counter$count = 82967;
	#10 counter$count = 82968;
	#10 counter$count = 82969;
	#10 counter$count = 82970;
	#10 counter$count = 82971;
	#10 counter$count = 82972;
	#10 counter$count = 82973;
	#10 counter$count = 82974;
	#10 counter$count = 82975;
	#10 counter$count = 82976;
	#10 counter$count = 82977;
	#10 counter$count = 82978;
	#10 counter$count = 82979;
	#10 counter$count = 82980;
	#10 counter$count = 82981;
	#10 counter$count = 82982;
	#10 counter$count = 82983;
	#10 counter$count = 82984;
	#10 counter$count = 82985;
	#10 counter$count = 82986;
	#10 counter$count = 82987;
	#10 counter$count = 82988;
	#10 counter$count = 82989;
	#10 counter$count = 82990;
	#10 counter$count = 82991;
	#10 counter$count = 82992;
	#10 counter$count = 82993;
	#10 counter$count = 82994;
	#10 counter$count = 82995;
	#10 counter$count = 82996;
	#10 counter$count = 82997;
	#10 counter$count = 82998;
	#10 counter$count = 82999;
	#10 counter$count = 83000;
	#10 counter$count = 83001;
	#10 counter$count = 83002;
	#10 counter$count = 83003;
	#10 counter$count = 83004;
	#10 counter$count = 83005;
	#10 counter$count = 83006;
	#10 counter$count = 83007;
	#10 counter$count = 83008;
	#10 counter$count = 83009;
	#10 counter$count = 83010;
	#10 counter$count = 83011;
	#10 counter$count = 83012;
	#10 counter$count = 83013;
	#10 counter$count = 83014;
	#10 counter$count = 83015;
	#10 counter$count = 83016;
	#10 counter$count = 83017;
	#10 counter$count = 83018;
	#10 counter$count = 83019;
	#10 counter$count = 83020;
	#10 counter$count = 83021;
	#10 counter$count = 83022;
	#10 counter$count = 83023;
	#10 counter$count = 83024;
	#10 counter$count = 83025;
	#10 counter$count = 83026;
	#10 counter$count = 83027;
	#10 counter$count = 83028;
	#10 counter$count = 83029;
	#10 counter$count = 83030;
	#10 counter$count = 83031;
	#10 counter$count = 83032;
	#10 counter$count = 83033;
	#10 counter$count = 83034;
	#10 counter$count = 83035;
	#10 counter$count = 83036;
	#10 counter$count = 83037;
	#10 counter$count = 83038;
	#10 counter$count = 83039;
	#10 counter$count = 83040;
	#10 counter$count = 83041;
	#10 counter$count = 83042;
	#10 counter$count = 83043;
	#10 counter$count = 83044;
	#10 counter$count = 83045;
	#10 counter$count = 83046;
	#10 counter$count = 83047;
	#10 counter$count = 83048;
	#10 counter$count = 83049;
	#10 counter$count = 83050;
	#10 counter$count = 83051;
	#10 counter$count = 83052;
	#10 counter$count = 83053;
	#10 counter$count = 83054;
	#10 counter$count = 83055;
	#10 counter$count = 83056;
	#10 counter$count = 83057;
	#10 counter$count = 83058;
	#10 counter$count = 83059;
	#10 counter$count = 83060;
	#10 counter$count = 83061;
	#10 counter$count = 83062;
	#10 counter$count = 83063;
	#10 counter$count = 83064;
	#10 counter$count = 83065;
	#10 counter$count = 83066;
	#10 counter$count = 83067;
	#10 counter$count = 83068;
	#10 counter$count = 83069;
	#10 counter$count = 83070;
	#10 counter$count = 83071;
	#10 counter$count = 83072;
	#10 counter$count = 83073;
	#10 counter$count = 83074;
	#10 counter$count = 83075;
	#10 counter$count = 83076;
	#10 counter$count = 83077;
	#10 counter$count = 83078;
	#10 counter$count = 83079;
	#10 counter$count = 83080;
	#10 counter$count = 83081;
	#10 counter$count = 83082;
	#10 counter$count = 83083;
	#10 counter$count = 83084;
	#10 counter$count = 83085;
	#10 counter$count = 83086;
	#10 counter$count = 83087;
	#10 counter$count = 83088;
	#10 counter$count = 83089;
	#10 counter$count = 83090;
	#10 counter$count = 83091;
	#10 counter$count = 83092;
	#10 counter$count = 83093;
	#10 counter$count = 83094;
	#10 counter$count = 83095;
	#10 counter$count = 83096;
	#10 counter$count = 83097;
	#10 counter$count = 83098;
	#10 counter$count = 83099;
	#10 counter$count = 83100;
	#10 counter$count = 83101;
	#10 counter$count = 83102;
	#10 counter$count = 83103;
	#10 counter$count = 83104;
	#10 counter$count = 83105;
	#10 counter$count = 83106;
	#10 counter$count = 83107;
	#10 counter$count = 83108;
	#10 counter$count = 83109;
	#10 counter$count = 83110;
	#10 counter$count = 83111;
	#10 counter$count = 83112;
	#10 counter$count = 83113;
	#10 counter$count = 83114;
	#10 counter$count = 83115;
	#10 counter$count = 83116;
	#10 counter$count = 83117;
	#10 counter$count = 83118;
	#10 counter$count = 83119;
	#10 counter$count = 83120;
	#10 counter$count = 83121;
	#10 counter$count = 83122;
	#10 counter$count = 83123;
	#10 counter$count = 83124;
	#10 counter$count = 83125;
	#10 counter$count = 83126;
	#10 counter$count = 83127;
	#10 counter$count = 83128;
	#10 counter$count = 83129;
	#10 counter$count = 83130;
	#10 counter$count = 83131;
	#10 counter$count = 83132;
	#10 counter$count = 83133;
	#10 counter$count = 83134;
	#10 counter$count = 83135;
	#10 counter$count = 83136;
	#10 counter$count = 83137;
	#10 counter$count = 83138;
	#10 counter$count = 83139;
	#10 counter$count = 83140;
	#10 counter$count = 83141;
	#10 counter$count = 83142;
	#10 counter$count = 83143;
	#10 counter$count = 83144;
	#10 counter$count = 83145;
	#10 counter$count = 83146;
	#10 counter$count = 83147;
	#10 counter$count = 83148;
	#10 counter$count = 83149;
	#10 counter$count = 83150;
	#10 counter$count = 83151;
	#10 counter$count = 83152;
	#10 counter$count = 83153;
	#10 counter$count = 83154;
	#10 counter$count = 83155;
	#10 counter$count = 83156;
	#10 counter$count = 83157;
	#10 counter$count = 83158;
	#10 counter$count = 83159;
	#10 counter$count = 83160;
	#10 counter$count = 83161;
	#10 counter$count = 83162;
	#10 counter$count = 83163;
	#10 counter$count = 83164;
	#10 counter$count = 83165;
	#10 counter$count = 83166;
	#10 counter$count = 83167;
	#10 counter$count = 83168;
	#10 counter$count = 83169;
	#10 counter$count = 83170;
	#10 counter$count = 83171;
	#10 counter$count = 83172;
	#10 counter$count = 83173;
	#10 counter$count = 83174;
	#10 counter$count = 83175;
	#10 counter$count = 83176;
	#10 counter$count = 83177;
	#10 counter$count = 83178;
	#10 counter$count = 83179;
	#10 counter$count = 83180;
	#10 counter$count = 83181;
	#10 counter$count = 83182;
	#10 counter$count = 83183;
	#10 counter$count = 83184;
	#10 counter$count = 83185;
	#10 counter$count = 83186;
	#10 counter$count = 83187;
	#10 counter$count = 83188;
	#10 counter$count = 83189;
	#10 counter$count = 83190;
	#10 counter$count = 83191;
	#10 counter$count = 83192;
	#10 counter$count = 83193;
	#10 counter$count = 83194;
	#10 counter$count = 83195;
	#10 counter$count = 83196;
	#10 counter$count = 83197;
	#10 counter$count = 83198;
	#10 counter$count = 83199;
	#10 counter$count = 83200;
	#10 counter$count = 83201;
	#10 counter$count = 83202;
	#10 counter$count = 83203;
	#10 counter$count = 83204;
	#10 counter$count = 83205;
	#10 counter$count = 83206;
	#10 counter$count = 83207;
	#10 counter$count = 83208;
	#10 counter$count = 83209;
	#10 counter$count = 83210;
	#10 counter$count = 83211;
	#10 counter$count = 83212;
	#10 counter$count = 83213;
	#10 counter$count = 83214;
	#10 counter$count = 83215;
	#10 counter$count = 83216;
	#10 counter$count = 83217;
	#10 counter$count = 83218;
	#10 counter$count = 83219;
	#10 counter$count = 83220;
	#10 counter$count = 83221;
	#10 counter$count = 83222;
	#10 counter$count = 83223;
	#10 counter$count = 83224;
	#10 counter$count = 83225;
	#10 counter$count = 83226;
	#10 counter$count = 83227;
	#10 counter$count = 83228;
	#10 counter$count = 83229;
	#10 counter$count = 83230;
	#10 counter$count = 83231;
	#10 counter$count = 83232;
	#10 counter$count = 83233;
	#10 counter$count = 83234;
	#10 counter$count = 83235;
	#10 counter$count = 83236;
	#10 counter$count = 83237;
	#10 counter$count = 83238;
	#10 counter$count = 83239;
	#10 counter$count = 83240;
	#10 counter$count = 83241;
	#10 counter$count = 83242;
	#10 counter$count = 83243;
	#10 counter$count = 83244;
	#10 counter$count = 83245;
	#10 counter$count = 83246;
	#10 counter$count = 83247;
	#10 counter$count = 83248;
	#10 counter$count = 83249;
	#10 counter$count = 83250;
	#10 counter$count = 83251;
	#10 counter$count = 83252;
	#10 counter$count = 83253;
	#10 counter$count = 83254;
	#10 counter$count = 83255;
	#10 counter$count = 83256;
	#10 counter$count = 83257;
	#10 counter$count = 83258;
	#10 counter$count = 83259;
	#10 counter$count = 83260;
	#10 counter$count = 83261;
	#10 counter$count = 83262;
	#10 counter$count = 83263;
	#10 counter$count = 83264;
	#10 counter$count = 83265;
	#10 counter$count = 83266;
	#10 counter$count = 83267;
	#10 counter$count = 83268;
	#10 counter$count = 83269;
	#10 counter$count = 83270;
	#10 counter$count = 83271;
	#10 counter$count = 83272;
	#10 counter$count = 83273;
	#10 counter$count = 83274;
	#10 counter$count = 83275;
	#10 counter$count = 83276;
	#10 counter$count = 83277;
	#10 counter$count = 83278;
	#10 counter$count = 83279;
	#10 counter$count = 83280;
	#10 counter$count = 83281;
	#10 counter$count = 83282;
	#10 counter$count = 83283;
	#10 counter$count = 83284;
	#10 counter$count = 83285;
	#10 counter$count = 83286;
	#10 counter$count = 83287;
	#10 counter$count = 83288;
	#10 counter$count = 83289;
	#10 counter$count = 83290;
	#10 counter$count = 83291;
	#10 counter$count = 83292;
	#10 counter$count = 83293;
	#10 counter$count = 83294;
	#10 counter$count = 83295;
	#10 counter$count = 83296;
	#10 counter$count = 83297;
	#10 counter$count = 83298;
	#10 counter$count = 83299;
	#10 counter$count = 83300;
	#10 counter$count = 83301;
	#10 counter$count = 83302;
	#10 counter$count = 83303;
	#10 counter$count = 83304;
	#10 counter$count = 83305;
	#10 counter$count = 83306;
	#10 counter$count = 83307;
	#10 counter$count = 83308;
	#10 counter$count = 83309;
	#10 counter$count = 83310;
	#10 counter$count = 83311;
	#10 counter$count = 83312;
	#10 counter$count = 83313;
	#10 counter$count = 83314;
	#10 counter$count = 83315;
	#10 counter$count = 83316;
	#10 counter$count = 83317;
	#10 counter$count = 83318;
	#10 counter$count = 83319;
	#10 counter$count = 83320;
	#10 counter$count = 83321;
	#10 counter$count = 83322;
	#10 counter$count = 83323;
	#10 counter$count = 83324;
	#10 counter$count = 83325;
	#10 counter$count = 83326;
	#10 counter$count = 83327;
	#10 counter$count = 83328;
	#10 counter$count = 83329;
	#10 counter$count = 83330;
	#10 counter$count = 83331;
	#10 counter$count = 83332;
	#10 counter$count = 83333;
	#10 counter$count = 83334;
	#10 counter$count = 83335;
	#10 counter$count = 83336;
	#10 counter$count = 83337;
	#10 counter$count = 83338;
	#10 counter$count = 83339;
	#10 counter$count = 83340;
	#10 counter$count = 83341;
	#10 counter$count = 83342;
	#10 counter$count = 83343;
	#10 counter$count = 83344;
	#10 counter$count = 83345;
	#10 counter$count = 83346;
	#10 counter$count = 83347;
	#10 counter$count = 83348;
	#10 counter$count = 83349;
	#10 counter$count = 83350;
	#10 counter$count = 83351;
	#10 counter$count = 83352;
	#10 counter$count = 83353;
	#10 counter$count = 83354;
	#10 counter$count = 83355;
	#10 counter$count = 83356;
	#10 counter$count = 83357;
	#10 counter$count = 83358;
	#10 counter$count = 83359;
	#10 counter$count = 83360;
	#10 counter$count = 83361;
	#10 counter$count = 83362;
	#10 counter$count = 83363;
	#10 counter$count = 83364;
	#10 counter$count = 83365;
	#10 counter$count = 83366;
	#10 counter$count = 83367;
	#10 counter$count = 83368;
	#10 counter$count = 83369;
	#10 counter$count = 83370;
	#10 counter$count = 83371;
	#10 counter$count = 83372;
	#10 counter$count = 83373;
	#10 counter$count = 83374;
	#10 counter$count = 83375;
	#10 counter$count = 83376;
	#10 counter$count = 83377;
	#10 counter$count = 83378;
	#10 counter$count = 83379;
	#10 counter$count = 83380;
	#10 counter$count = 83381;
	#10 counter$count = 83382;
	#10 counter$count = 83383;
	#10 counter$count = 83384;
	#10 counter$count = 83385;
	#10 counter$count = 83386;
	#10 counter$count = 83387;
	#10 counter$count = 83388;
	#10 counter$count = 83389;
	#10 counter$count = 83390;
	#10 counter$count = 83391;
	#10 counter$count = 83392;
	#10 counter$count = 83393;
	#10 counter$count = 83394;
	#10 counter$count = 83395;
	#10 counter$count = 83396;
	#10 counter$count = 83397;
	#10 counter$count = 83398;
	#10 counter$count = 83399;
	#10 counter$count = 83400;
	#10 counter$count = 83401;
	#10 counter$count = 83402;
	#10 counter$count = 83403;
	#10 counter$count = 83404;
	#10 counter$count = 83405;
	#10 counter$count = 83406;
	#10 counter$count = 83407;
	#10 counter$count = 83408;
	#10 counter$count = 83409;
	#10 counter$count = 83410;
	#10 counter$count = 83411;
	#10 counter$count = 83412;
	#10 counter$count = 83413;
	#10 counter$count = 83414;
	#10 counter$count = 83415;
	#10 counter$count = 83416;
	#10 counter$count = 83417;
	#10 counter$count = 83418;
	#10 counter$count = 83419;
	#10 counter$count = 83420;
	#10 counter$count = 83421;
	#10 counter$count = 83422;
	#10 counter$count = 83423;
	#10 counter$count = 83424;
	#10 counter$count = 83425;
	#10 counter$count = 83426;
	#10 counter$count = 83427;
	#10 counter$count = 83428;
	#10 counter$count = 83429;
	#10 counter$count = 83430;
	#10 counter$count = 83431;
	#10 counter$count = 83432;
	#10 counter$count = 83433;
	#10 counter$count = 83434;
	#10 counter$count = 83435;
	#10 counter$count = 83436;
	#10 counter$count = 83437;
	#10 counter$count = 83438;
	#10 counter$count = 83439;
	#10 counter$count = 83440;
	#10 counter$count = 83441;
	#10 counter$count = 83442;
	#10 counter$count = 83443;
	#10 counter$count = 83444;
	#10 counter$count = 83445;
	#10 counter$count = 83446;
	#10 counter$count = 83447;
	#10 counter$count = 83448;
	#10 counter$count = 83449;
	#10 counter$count = 83450;
	#10 counter$count = 83451;
	#10 counter$count = 83452;
	#10 counter$count = 83453;
	#10 counter$count = 83454;
	#10 counter$count = 83455;
	#10 counter$count = 83456;
	#10 counter$count = 83457;
	#10 counter$count = 83458;
	#10 counter$count = 83459;
	#10 counter$count = 83460;
	#10 counter$count = 83461;
	#10 counter$count = 83462;
	#10 counter$count = 83463;
	#10 counter$count = 83464;
	#10 counter$count = 83465;
	#10 counter$count = 83466;
	#10 counter$count = 83467;
	#10 counter$count = 83468;
	#10 counter$count = 83469;
	#10 counter$count = 83470;
	#10 counter$count = 83471;
	#10 counter$count = 83472;
	#10 counter$count = 83473;
	#10 counter$count = 83474;
	#10 counter$count = 83475;
	#10 counter$count = 83476;
	#10 counter$count = 83477;
	#10 counter$count = 83478;
	#10 counter$count = 83479;
	#10 counter$count = 83480;
	#10 counter$count = 83481;
	#10 counter$count = 83482;
	#10 counter$count = 83483;
	#10 counter$count = 83484;
	#10 counter$count = 83485;
	#10 counter$count = 83486;
	#10 counter$count = 83487;
	#10 counter$count = 83488;
	#10 counter$count = 83489;
	#10 counter$count = 83490;
	#10 counter$count = 83491;
	#10 counter$count = 83492;
	#10 counter$count = 83493;
	#10 counter$count = 83494;
	#10 counter$count = 83495;
	#10 counter$count = 83496;
	#10 counter$count = 83497;
	#10 counter$count = 83498;
	#10 counter$count = 83499;
	#10 counter$count = 83500;
	#10 counter$count = 83501;
	#10 counter$count = 83502;
	#10 counter$count = 83503;
	#10 counter$count = 83504;
	#10 counter$count = 83505;
	#10 counter$count = 83506;
	#10 counter$count = 83507;
	#10 counter$count = 83508;
	#10 counter$count = 83509;
	#10 counter$count = 83510;
	#10 counter$count = 83511;
	#10 counter$count = 83512;
	#10 counter$count = 83513;
	#10 counter$count = 83514;
	#10 counter$count = 83515;
	#10 counter$count = 83516;
	#10 counter$count = 83517;
	#10 counter$count = 83518;
	#10 counter$count = 83519;
	#10 counter$count = 83520;
	#10 counter$count = 83521;
	#10 counter$count = 83522;
	#10 counter$count = 83523;
	#10 counter$count = 83524;
	#10 counter$count = 83525;
	#10 counter$count = 83526;
	#10 counter$count = 83527;
	#10 counter$count = 83528;
	#10 counter$count = 83529;
	#10 counter$count = 83530;
	#10 counter$count = 83531;
	#10 counter$count = 83532;
	#10 counter$count = 83533;
	#10 counter$count = 83534;
	#10 counter$count = 83535;
	#10 counter$count = 83536;
	#10 counter$count = 83537;
	#10 counter$count = 83538;
	#10 counter$count = 83539;
	#10 counter$count = 83540;
	#10 counter$count = 83541;
	#10 counter$count = 83542;
	#10 counter$count = 83543;
	#10 counter$count = 83544;
	#10 counter$count = 83545;
	#10 counter$count = 83546;
	#10 counter$count = 83547;
	#10 counter$count = 83548;
	#10 counter$count = 83549;
	#10 counter$count = 83550;
	#10 counter$count = 83551;
	#10 counter$count = 83552;
	#10 counter$count = 83553;
	#10 counter$count = 83554;
	#10 counter$count = 83555;
	#10 counter$count = 83556;
	#10 counter$count = 83557;
	#10 counter$count = 83558;
	#10 counter$count = 83559;
	#10 counter$count = 83560;
	#10 counter$count = 83561;
	#10 counter$count = 83562;
	#10 counter$count = 83563;
	#10 counter$count = 83564;
	#10 counter$count = 83565;
	#10 counter$count = 83566;
	#10 counter$count = 83567;
	#10 counter$count = 83568;
	#10 counter$count = 83569;
	#10 counter$count = 83570;
	#10 counter$count = 83571;
	#10 counter$count = 83572;
	#10 counter$count = 83573;
	#10 counter$count = 83574;
	#10 counter$count = 83575;
	#10 counter$count = 83576;
	#10 counter$count = 83577;
	#10 counter$count = 83578;
	#10 counter$count = 83579;
	#10 counter$count = 83580;
	#10 counter$count = 83581;
	#10 counter$count = 83582;
	#10 counter$count = 83583;
	#10 counter$count = 83584;
	#10 counter$count = 83585;
	#10 counter$count = 83586;
	#10 counter$count = 83587;
	#10 counter$count = 83588;
	#10 counter$count = 83589;
	#10 counter$count = 83590;
	#10 counter$count = 83591;
	#10 counter$count = 83592;
	#10 counter$count = 83593;
	#10 counter$count = 83594;
	#10 counter$count = 83595;
	#10 counter$count = 83596;
	#10 counter$count = 83597;
	#10 counter$count = 83598;
	#10 counter$count = 83599;
	#10 counter$count = 83600;
	#10 counter$count = 83601;
	#10 counter$count = 83602;
	#10 counter$count = 83603;
	#10 counter$count = 83604;
	#10 counter$count = 83605;
	#10 counter$count = 83606;
	#10 counter$count = 83607;
	#10 counter$count = 83608;
	#10 counter$count = 83609;
	#10 counter$count = 83610;
	#10 counter$count = 83611;
	#10 counter$count = 83612;
	#10 counter$count = 83613;
	#10 counter$count = 83614;
	#10 counter$count = 83615;
	#10 counter$count = 83616;
	#10 counter$count = 83617;
	#10 counter$count = 83618;
	#10 counter$count = 83619;
	#10 counter$count = 83620;
	#10 counter$count = 83621;
	#10 counter$count = 83622;
	#10 counter$count = 83623;
	#10 counter$count = 83624;
	#10 counter$count = 83625;
	#10 counter$count = 83626;
	#10 counter$count = 83627;
	#10 counter$count = 83628;
	#10 counter$count = 83629;
	#10 counter$count = 83630;
	#10 counter$count = 83631;
	#10 counter$count = 83632;
	#10 counter$count = 83633;
	#10 counter$count = 83634;
	#10 counter$count = 83635;
	#10 counter$count = 83636;
	#10 counter$count = 83637;
	#10 counter$count = 83638;
	#10 counter$count = 83639;
	#10 counter$count = 83640;
	#10 counter$count = 83641;
	#10 counter$count = 83642;
	#10 counter$count = 83643;
	#10 counter$count = 83644;
	#10 counter$count = 83645;
	#10 counter$count = 83646;
	#10 counter$count = 83647;
	#10 counter$count = 83648;
	#10 counter$count = 83649;
	#10 counter$count = 83650;
	#10 counter$count = 83651;
	#10 counter$count = 83652;
	#10 counter$count = 83653;
	#10 counter$count = 83654;
	#10 counter$count = 83655;
	#10 counter$count = 83656;
	#10 counter$count = 83657;
	#10 counter$count = 83658;
	#10 counter$count = 83659;
	#10 counter$count = 83660;
	#10 counter$count = 83661;
	#10 counter$count = 83662;
	#10 counter$count = 83663;
	#10 counter$count = 83664;
	#10 counter$count = 83665;
	#10 counter$count = 83666;
	#10 counter$count = 83667;
	#10 counter$count = 83668;
	#10 counter$count = 83669;
	#10 counter$count = 83670;
	#10 counter$count = 83671;
	#10 counter$count = 83672;
	#10 counter$count = 83673;
	#10 counter$count = 83674;
	#10 counter$count = 83675;
	#10 counter$count = 83676;
	#10 counter$count = 83677;
	#10 counter$count = 83678;
	#10 counter$count = 83679;
	#10 counter$count = 83680;
	#10 counter$count = 83681;
	#10 counter$count = 83682;
	#10 counter$count = 83683;
	#10 counter$count = 83684;
	#10 counter$count = 83685;
	#10 counter$count = 83686;
	#10 counter$count = 83687;
	#10 counter$count = 83688;
	#10 counter$count = 83689;
	#10 counter$count = 83690;
	#10 counter$count = 83691;
	#10 counter$count = 83692;
	#10 counter$count = 83693;
	#10 counter$count = 83694;
	#10 counter$count = 83695;
	#10 counter$count = 83696;
	#10 counter$count = 83697;
	#10 counter$count = 83698;
	#10 counter$count = 83699;
	#10 counter$count = 83700;
	#10 counter$count = 83701;
	#10 counter$count = 83702;
	#10 counter$count = 83703;
	#10 counter$count = 83704;
	#10 counter$count = 83705;
	#10 counter$count = 83706;
	#10 counter$count = 83707;
	#10 counter$count = 83708;
	#10 counter$count = 83709;
	#10 counter$count = 83710;
	#10 counter$count = 83711;
	#10 counter$count = 83712;
	#10 counter$count = 83713;
	#10 counter$count = 83714;
	#10 counter$count = 83715;
	#10 counter$count = 83716;
	#10 counter$count = 83717;
	#10 counter$count = 83718;
	#10 counter$count = 83719;
	#10 counter$count = 83720;
	#10 counter$count = 83721;
	#10 counter$count = 83722;
	#10 counter$count = 83723;
	#10 counter$count = 83724;
	#10 counter$count = 83725;
	#10 counter$count = 83726;
	#10 counter$count = 83727;
	#10 counter$count = 83728;
	#10 counter$count = 83729;
	#10 counter$count = 83730;
	#10 counter$count = 83731;
	#10 counter$count = 83732;
	#10 counter$count = 83733;
	#10 counter$count = 83734;
	#10 counter$count = 83735;
	#10 counter$count = 83736;
	#10 counter$count = 83737;
	#10 counter$count = 83738;
	#10 counter$count = 83739;
	#10 counter$count = 83740;
	#10 counter$count = 83741;
	#10 counter$count = 83742;
	#10 counter$count = 83743;
	#10 counter$count = 83744;
	#10 counter$count = 83745;
	#10 counter$count = 83746;
	#10 counter$count = 83747;
	#10 counter$count = 83748;
	#10 counter$count = 83749;
	#10 counter$count = 83750;
	#10 counter$count = 83751;
	#10 counter$count = 83752;
	#10 counter$count = 83753;
	#10 counter$count = 83754;
	#10 counter$count = 83755;
	#10 counter$count = 83756;
	#10 counter$count = 83757;
	#10 counter$count = 83758;
	#10 counter$count = 83759;
	#10 counter$count = 83760;
	#10 counter$count = 83761;
	#10 counter$count = 83762;
	#10 counter$count = 83763;
	#10 counter$count = 83764;
	#10 counter$count = 83765;
	#10 counter$count = 83766;
	#10 counter$count = 83767;
	#10 counter$count = 83768;
	#10 counter$count = 83769;
	#10 counter$count = 83770;
	#10 counter$count = 83771;
	#10 counter$count = 83772;
	#10 counter$count = 83773;
	#10 counter$count = 83774;
	#10 counter$count = 83775;
	#10 counter$count = 83776;
	#10 counter$count = 83777;
	#10 counter$count = 83778;
	#10 counter$count = 83779;
	#10 counter$count = 83780;
	#10 counter$count = 83781;
	#10 counter$count = 83782;
	#10 counter$count = 83783;
	#10 counter$count = 83784;
	#10 counter$count = 83785;
	#10 counter$count = 83786;
	#10 counter$count = 83787;
	#10 counter$count = 83788;
	#10 counter$count = 83789;
	#10 counter$count = 83790;
	#10 counter$count = 83791;
	#10 counter$count = 83792;
	#10 counter$count = 83793;
	#10 counter$count = 83794;
	#10 counter$count = 83795;
	#10 counter$count = 83796;
	#10 counter$count = 83797;
	#10 counter$count = 83798;
	#10 counter$count = 83799;
	#10 counter$count = 83800;
	#10 counter$count = 83801;
	#10 counter$count = 83802;
	#10 counter$count = 83803;
	#10 counter$count = 83804;
	#10 counter$count = 83805;
	#10 counter$count = 83806;
	#10 counter$count = 83807;
	#10 counter$count = 83808;
	#10 counter$count = 83809;
	#10 counter$count = 83810;
	#10 counter$count = 83811;
	#10 counter$count = 83812;
	#10 counter$count = 83813;
	#10 counter$count = 83814;
	#10 counter$count = 83815;
	#10 counter$count = 83816;
	#10 counter$count = 83817;
	#10 counter$count = 83818;
	#10 counter$count = 83819;
	#10 counter$count = 83820;
	#10 counter$count = 83821;
	#10 counter$count = 83822;
	#10 counter$count = 83823;
	#10 counter$count = 83824;
	#10 counter$count = 83825;
	#10 counter$count = 83826;
	#10 counter$count = 83827;
	#10 counter$count = 83828;
	#10 counter$count = 83829;
	#10 counter$count = 83830;
	#10 counter$count = 83831;
	#10 counter$count = 83832;
	#10 counter$count = 83833;
	#10 counter$count = 83834;
	#10 counter$count = 83835;
	#10 counter$count = 83836;
	#10 counter$count = 83837;
	#10 counter$count = 83838;
	#10 counter$count = 83839;
	#10 counter$count = 83840;
	#10 counter$count = 83841;
	#10 counter$count = 83842;
	#10 counter$count = 83843;
	#10 counter$count = 83844;
	#10 counter$count = 83845;
	#10 counter$count = 83846;
	#10 counter$count = 83847;
	#10 counter$count = 83848;
	#10 counter$count = 83849;
	#10 counter$count = 83850;
	#10 counter$count = 83851;
	#10 counter$count = 83852;
	#10 counter$count = 83853;
	#10 counter$count = 83854;
	#10 counter$count = 83855;
	#10 counter$count = 83856;
	#10 counter$count = 83857;
	#10 counter$count = 83858;
	#10 counter$count = 83859;
	#10 counter$count = 83860;
	#10 counter$count = 83861;
	#10 counter$count = 83862;
	#10 counter$count = 83863;
	#10 counter$count = 83864;
	#10 counter$count = 83865;
	#10 counter$count = 83866;
	#10 counter$count = 83867;
	#10 counter$count = 83868;
	#10 counter$count = 83869;
	#10 counter$count = 83870;
	#10 counter$count = 83871;
	#10 counter$count = 83872;
	#10 counter$count = 83873;
	#10 counter$count = 83874;
	#10 counter$count = 83875;
	#10 counter$count = 83876;
	#10 counter$count = 83877;
	#10 counter$count = 83878;
	#10 counter$count = 83879;
	#10 counter$count = 83880;
	#10 counter$count = 83881;
	#10 counter$count = 83882;
	#10 counter$count = 83883;
	#10 counter$count = 83884;
	#10 counter$count = 83885;
	#10 counter$count = 83886;
	#10 counter$count = 83887;
	#10 counter$count = 83888;
	#10 counter$count = 83889;
	#10 counter$count = 83890;
	#10 counter$count = 83891;
	#10 counter$count = 83892;
	#10 counter$count = 83893;
	#10 counter$count = 83894;
	#10 counter$count = 83895;
	#10 counter$count = 83896;
	#10 counter$count = 83897;
	#10 counter$count = 83898;
	#10 counter$count = 83899;
	#10 counter$count = 83900;
	#10 counter$count = 83901;
	#10 counter$count = 83902;
	#10 counter$count = 83903;
	#10 counter$count = 83904;
	#10 counter$count = 83905;
	#10 counter$count = 83906;
	#10 counter$count = 83907;
	#10 counter$count = 83908;
	#10 counter$count = 83909;
	#10 counter$count = 83910;
	#10 counter$count = 83911;
	#10 counter$count = 83912;
	#10 counter$count = 83913;
	#10 counter$count = 83914;
	#10 counter$count = 83915;
	#10 counter$count = 83916;
	#10 counter$count = 83917;
	#10 counter$count = 83918;
	#10 counter$count = 83919;
	#10 counter$count = 83920;
	#10 counter$count = 83921;
	#10 counter$count = 83922;
	#10 counter$count = 83923;
	#10 counter$count = 83924;
	#10 counter$count = 83925;
	#10 counter$count = 83926;
	#10 counter$count = 83927;
	#10 counter$count = 83928;
	#10 counter$count = 83929;
	#10 counter$count = 83930;
	#10 counter$count = 83931;
	#10 counter$count = 83932;
	#10 counter$count = 83933;
	#10 counter$count = 83934;
	#10 counter$count = 83935;
	#10 counter$count = 83936;
	#10 counter$count = 83937;
	#10 counter$count = 83938;
	#10 counter$count = 83939;
	#10 counter$count = 83940;
	#10 counter$count = 83941;
	#10 counter$count = 83942;
	#10 counter$count = 83943;
	#10 counter$count = 83944;
	#10 counter$count = 83945;
	#10 counter$count = 83946;
	#10 counter$count = 83947;
	#10 counter$count = 83948;
	#10 counter$count = 83949;
	#10 counter$count = 83950;
	#10 counter$count = 83951;
	#10 counter$count = 83952;
	#10 counter$count = 83953;
	#10 counter$count = 83954;
	#10 counter$count = 83955;
	#10 counter$count = 83956;
	#10 counter$count = 83957;
	#10 counter$count = 83958;
	#10 counter$count = 83959;
	#10 counter$count = 83960;
	#10 counter$count = 83961;
	#10 counter$count = 83962;
	#10 counter$count = 83963;
	#10 counter$count = 83964;
	#10 counter$count = 83965;
	#10 counter$count = 83966;
	#10 counter$count = 83967;
	#10 counter$count = 83968;
	#10 counter$count = 83969;
	#10 counter$count = 83970;
	#10 counter$count = 83971;
	#10 counter$count = 83972;
	#10 counter$count = 83973;
	#10 counter$count = 83974;
	#10 counter$count = 83975;
	#10 counter$count = 83976;
	#10 counter$count = 83977;
	#10 counter$count = 83978;
	#10 counter$count = 83979;
	#10 counter$count = 83980;
	#10 counter$count = 83981;
	#10 counter$count = 83982;
	#10 counter$count = 83983;
	#10 counter$count = 83984;
	#10 counter$count = 83985;
	#10 counter$count = 83986;
	#10 counter$count = 83987;
	#10 counter$count = 83988;
	#10 counter$count = 83989;
	#10 counter$count = 83990;
	#10 counter$count = 83991;
	#10 counter$count = 83992;
	#10 counter$count = 83993;
	#10 counter$count = 83994;
	#10 counter$count = 83995;
	#10 counter$count = 83996;
	#10 counter$count = 83997;
	#10 counter$count = 83998;
	#10 counter$count = 83999;
	#10 counter$count = 84000;
	#10 counter$count = 84001;
	#10 counter$count = 84002;
	#10 counter$count = 84003;
	#10 counter$count = 84004;
	#10 counter$count = 84005;
	#10 counter$count = 84006;
	#10 counter$count = 84007;
	#10 counter$count = 84008;
	#10 counter$count = 84009;
	#10 counter$count = 84010;
	#10 counter$count = 84011;
	#10 counter$count = 84012;
	#10 counter$count = 84013;
	#10 counter$count = 84014;
	#10 counter$count = 84015;
	#10 counter$count = 84016;
	#10 counter$count = 84017;
	#10 counter$count = 84018;
	#10 counter$count = 84019;
	#10 counter$count = 84020;
	#10 counter$count = 84021;
	#10 counter$count = 84022;
	#10 counter$count = 84023;
	#10 counter$count = 84024;
	#10 counter$count = 84025;
	#10 counter$count = 84026;
	#10 counter$count = 84027;
	#10 counter$count = 84028;
	#10 counter$count = 84029;
	#10 counter$count = 84030;
	#10 counter$count = 84031;
	#10 counter$count = 84032;
	#10 counter$count = 84033;
	#10 counter$count = 84034;
	#10 counter$count = 84035;
	#10 counter$count = 84036;
	#10 counter$count = 84037;
	#10 counter$count = 84038;
	#10 counter$count = 84039;
	#10 counter$count = 84040;
	#10 counter$count = 84041;
	#10 counter$count = 84042;
	#10 counter$count = 84043;
	#10 counter$count = 84044;
	#10 counter$count = 84045;
	#10 counter$count = 84046;
	#10 counter$count = 84047;
	#10 counter$count = 84048;
	#10 counter$count = 84049;
	#10 counter$count = 84050;
	#10 counter$count = 84051;
	#10 counter$count = 84052;
	#10 counter$count = 84053;
	#10 counter$count = 84054;
	#10 counter$count = 84055;
	#10 counter$count = 84056;
	#10 counter$count = 84057;
	#10 counter$count = 84058;
	#10 counter$count = 84059;
	#10 counter$count = 84060;
	#10 counter$count = 84061;
	#10 counter$count = 84062;
	#10 counter$count = 84063;
	#10 counter$count = 84064;
	#10 counter$count = 84065;
	#10 counter$count = 84066;
	#10 counter$count = 84067;
	#10 counter$count = 84068;
	#10 counter$count = 84069;
	#10 counter$count = 84070;
	#10 counter$count = 84071;
	#10 counter$count = 84072;
	#10 counter$count = 84073;
	#10 counter$count = 84074;
	#10 counter$count = 84075;
	#10 counter$count = 84076;
	#10 counter$count = 84077;
	#10 counter$count = 84078;
	#10 counter$count = 84079;
	#10 counter$count = 84080;
	#10 counter$count = 84081;
	#10 counter$count = 84082;
	#10 counter$count = 84083;
	#10 counter$count = 84084;
	#10 counter$count = 84085;
	#10 counter$count = 84086;
	#10 counter$count = 84087;
	#10 counter$count = 84088;
	#10 counter$count = 84089;
	#10 counter$count = 84090;
	#10 counter$count = 84091;
	#10 counter$count = 84092;
	#10 counter$count = 84093;
	#10 counter$count = 84094;
	#10 counter$count = 84095;
	#10 counter$count = 84096;
	#10 counter$count = 84097;
	#10 counter$count = 84098;
	#10 counter$count = 84099;
	#10 counter$count = 84100;
	#10 counter$count = 84101;
	#10 counter$count = 84102;
	#10 counter$count = 84103;
	#10 counter$count = 84104;
	#10 counter$count = 84105;
	#10 counter$count = 84106;
	#10 counter$count = 84107;
	#10 counter$count = 84108;
	#10 counter$count = 84109;
	#10 counter$count = 84110;
	#10 counter$count = 84111;
	#10 counter$count = 84112;
	#10 counter$count = 84113;
	#10 counter$count = 84114;
	#10 counter$count = 84115;
	#10 counter$count = 84116;
	#10 counter$count = 84117;
	#10 counter$count = 84118;
	#10 counter$count = 84119;
	#10 counter$count = 84120;
	#10 counter$count = 84121;
	#10 counter$count = 84122;
	#10 counter$count = 84123;
	#10 counter$count = 84124;
	#10 counter$count = 84125;
	#10 counter$count = 84126;
	#10 counter$count = 84127;
	#10 counter$count = 84128;
	#10 counter$count = 84129;
	#10 counter$count = 84130;
	#10 counter$count = 84131;
	#10 counter$count = 84132;
	#10 counter$count = 84133;
	#10 counter$count = 84134;
	#10 counter$count = 84135;
	#10 counter$count = 84136;
	#10 counter$count = 84137;
	#10 counter$count = 84138;
	#10 counter$count = 84139;
	#10 counter$count = 84140;
	#10 counter$count = 84141;
	#10 counter$count = 84142;
	#10 counter$count = 84143;
	#10 counter$count = 84144;
	#10 counter$count = 84145;
	#10 counter$count = 84146;
	#10 counter$count = 84147;
	#10 counter$count = 84148;
	#10 counter$count = 84149;
	#10 counter$count = 84150;
	#10 counter$count = 84151;
	#10 counter$count = 84152;
	#10 counter$count = 84153;
	#10 counter$count = 84154;
	#10 counter$count = 84155;
	#10 counter$count = 84156;
	#10 counter$count = 84157;
	#10 counter$count = 84158;
	#10 counter$count = 84159;
	#10 counter$count = 84160;
	#10 counter$count = 84161;
	#10 counter$count = 84162;
	#10 counter$count = 84163;
	#10 counter$count = 84164;
	#10 counter$count = 84165;
	#10 counter$count = 84166;
	#10 counter$count = 84167;
	#10 counter$count = 84168;
	#10 counter$count = 84169;
	#10 counter$count = 84170;
	#10 counter$count = 84171;
	#10 counter$count = 84172;
	#10 counter$count = 84173;
	#10 counter$count = 84174;
	#10 counter$count = 84175;
	#10 counter$count = 84176;
	#10 counter$count = 84177;
	#10 counter$count = 84178;
	#10 counter$count = 84179;
	#10 counter$count = 84180;
	#10 counter$count = 84181;
	#10 counter$count = 84182;
	#10 counter$count = 84183;
	#10 counter$count = 84184;
	#10 counter$count = 84185;
	#10 counter$count = 84186;
	#10 counter$count = 84187;
	#10 counter$count = 84188;
	#10 counter$count = 84189;
	#10 counter$count = 84190;
	#10 counter$count = 84191;
	#10 counter$count = 84192;
	#10 counter$count = 84193;
	#10 counter$count = 84194;
	#10 counter$count = 84195;
	#10 counter$count = 84196;
	#10 counter$count = 84197;
	#10 counter$count = 84198;
	#10 counter$count = 84199;
	#10 counter$count = 84200;
	#10 counter$count = 84201;
	#10 counter$count = 84202;
	#10 counter$count = 84203;
	#10 counter$count = 84204;
	#10 counter$count = 84205;
	#10 counter$count = 84206;
	#10 counter$count = 84207;
	#10 counter$count = 84208;
	#10 counter$count = 84209;
	#10 counter$count = 84210;
	#10 counter$count = 84211;
	#10 counter$count = 84212;
	#10 counter$count = 84213;
	#10 counter$count = 84214;
	#10 counter$count = 84215;
	#10 counter$count = 84216;
	#10 counter$count = 84217;
	#10 counter$count = 84218;
	#10 counter$count = 84219;
	#10 counter$count = 84220;
	#10 counter$count = 84221;
	#10 counter$count = 84222;
	#10 counter$count = 84223;
	#10 counter$count = 84224;
	#10 counter$count = 84225;
	#10 counter$count = 84226;
	#10 counter$count = 84227;
	#10 counter$count = 84228;
	#10 counter$count = 84229;
	#10 counter$count = 84230;
	#10 counter$count = 84231;
	#10 counter$count = 84232;
	#10 counter$count = 84233;
	#10 counter$count = 84234;
	#10 counter$count = 84235;
	#10 counter$count = 84236;
	#10 counter$count = 84237;
	#10 counter$count = 84238;
	#10 counter$count = 84239;
	#10 counter$count = 84240;
	#10 counter$count = 84241;
	#10 counter$count = 84242;
	#10 counter$count = 84243;
	#10 counter$count = 84244;
	#10 counter$count = 84245;
	#10 counter$count = 84246;
	#10 counter$count = 84247;
	#10 counter$count = 84248;
	#10 counter$count = 84249;
	#10 counter$count = 84250;
	#10 counter$count = 84251;
	#10 counter$count = 84252;
	#10 counter$count = 84253;
	#10 counter$count = 84254;
	#10 counter$count = 84255;
	#10 counter$count = 84256;
	#10 counter$count = 84257;
	#10 counter$count = 84258;
	#10 counter$count = 84259;
	#10 counter$count = 84260;
	#10 counter$count = 84261;
	#10 counter$count = 84262;
	#10 counter$count = 84263;
	#10 counter$count = 84264;
	#10 counter$count = 84265;
	#10 counter$count = 84266;
	#10 counter$count = 84267;
	#10 counter$count = 84268;
	#10 counter$count = 84269;
	#10 counter$count = 84270;
	#10 counter$count = 84271;
	#10 counter$count = 84272;
	#10 counter$count = 84273;
	#10 counter$count = 84274;
	#10 counter$count = 84275;
	#10 counter$count = 84276;
	#10 counter$count = 84277;
	#10 counter$count = 84278;
	#10 counter$count = 84279;
	#10 counter$count = 84280;
	#10 counter$count = 84281;
	#10 counter$count = 84282;
	#10 counter$count = 84283;
	#10 counter$count = 84284;
	#10 counter$count = 84285;
	#10 counter$count = 84286;
	#10 counter$count = 84287;
	#10 counter$count = 84288;
	#10 counter$count = 84289;
	#10 counter$count = 84290;
	#10 counter$count = 84291;
	#10 counter$count = 84292;
	#10 counter$count = 84293;
	#10 counter$count = 84294;
	#10 counter$count = 84295;
	#10 counter$count = 84296;
	#10 counter$count = 84297;
	#10 counter$count = 84298;
	#10 counter$count = 84299;
	#10 counter$count = 84300;
	#10 counter$count = 84301;
	#10 counter$count = 84302;
	#10 counter$count = 84303;
	#10 counter$count = 84304;
	#10 counter$count = 84305;
	#10 counter$count = 84306;
	#10 counter$count = 84307;
	#10 counter$count = 84308;
	#10 counter$count = 84309;
	#10 counter$count = 84310;
	#10 counter$count = 84311;
	#10 counter$count = 84312;
	#10 counter$count = 84313;
	#10 counter$count = 84314;
	#10 counter$count = 84315;
	#10 counter$count = 84316;
	#10 counter$count = 84317;
	#10 counter$count = 84318;
	#10 counter$count = 84319;
	#10 counter$count = 84320;
	#10 counter$count = 84321;
	#10 counter$count = 84322;
	#10 counter$count = 84323;
	#10 counter$count = 84324;
	#10 counter$count = 84325;
	#10 counter$count = 84326;
	#10 counter$count = 84327;
	#10 counter$count = 84328;
	#10 counter$count = 84329;
	#10 counter$count = 84330;
	#10 counter$count = 84331;
	#10 counter$count = 84332;
	#10 counter$count = 84333;
	#10 counter$count = 84334;
	#10 counter$count = 84335;
	#10 counter$count = 84336;
	#10 counter$count = 84337;
	#10 counter$count = 84338;
	#10 counter$count = 84339;
	#10 counter$count = 84340;
	#10 counter$count = 84341;
	#10 counter$count = 84342;
	#10 counter$count = 84343;
	#10 counter$count = 84344;
	#10 counter$count = 84345;
	#10 counter$count = 84346;
	#10 counter$count = 84347;
	#10 counter$count = 84348;
	#10 counter$count = 84349;
	#10 counter$count = 84350;
	#10 counter$count = 84351;
	#10 counter$count = 84352;
	#10 counter$count = 84353;
	#10 counter$count = 84354;
	#10 counter$count = 84355;
	#10 counter$count = 84356;
	#10 counter$count = 84357;
	#10 counter$count = 84358;
	#10 counter$count = 84359;
	#10 counter$count = 84360;
	#10 counter$count = 84361;
	#10 counter$count = 84362;
	#10 counter$count = 84363;
	#10 counter$count = 84364;
	#10 counter$count = 84365;
	#10 counter$count = 84366;
	#10 counter$count = 84367;
	#10 counter$count = 84368;
	#10 counter$count = 84369;
	#10 counter$count = 84370;
	#10 counter$count = 84371;
	#10 counter$count = 84372;
	#10 counter$count = 84373;
	#10 counter$count = 84374;
	#10 counter$count = 84375;
	#10 counter$count = 84376;
	#10 counter$count = 84377;
	#10 counter$count = 84378;
	#10 counter$count = 84379;
	#10 counter$count = 84380;
	#10 counter$count = 84381;
	#10 counter$count = 84382;
	#10 counter$count = 84383;
	#10 counter$count = 84384;
	#10 counter$count = 84385;
	#10 counter$count = 84386;
	#10 counter$count = 84387;
	#10 counter$count = 84388;
	#10 counter$count = 84389;
	#10 counter$count = 84390;
	#10 counter$count = 84391;
	#10 counter$count = 84392;
	#10 counter$count = 84393;
	#10 counter$count = 84394;
	#10 counter$count = 84395;
	#10 counter$count = 84396;
	#10 counter$count = 84397;
	#10 counter$count = 84398;
	#10 counter$count = 84399;
	#10 counter$count = 84400;
	#10 counter$count = 84401;
	#10 counter$count = 84402;
	#10 counter$count = 84403;
	#10 counter$count = 84404;
	#10 counter$count = 84405;
	#10 counter$count = 84406;
	#10 counter$count = 84407;
	#10 counter$count = 84408;
	#10 counter$count = 84409;
	#10 counter$count = 84410;
	#10 counter$count = 84411;
	#10 counter$count = 84412;
	#10 counter$count = 84413;
	#10 counter$count = 84414;
	#10 counter$count = 84415;
	#10 counter$count = 84416;
	#10 counter$count = 84417;
	#10 counter$count = 84418;
	#10 counter$count = 84419;
	#10 counter$count = 84420;
	#10 counter$count = 84421;
	#10 counter$count = 84422;
	#10 counter$count = 84423;
	#10 counter$count = 84424;
	#10 counter$count = 84425;
	#10 counter$count = 84426;
	#10 counter$count = 84427;
	#10 counter$count = 84428;
	#10 counter$count = 84429;
	#10 counter$count = 84430;
	#10 counter$count = 84431;
	#10 counter$count = 84432;
	#10 counter$count = 84433;
	#10 counter$count = 84434;
	#10 counter$count = 84435;
	#10 counter$count = 84436;
	#10 counter$count = 84437;
	#10 counter$count = 84438;
	#10 counter$count = 84439;
	#10 counter$count = 84440;
	#10 counter$count = 84441;
	#10 counter$count = 84442;
	#10 counter$count = 84443;
	#10 counter$count = 84444;
	#10 counter$count = 84445;
	#10 counter$count = 84446;
	#10 counter$count = 84447;
	#10 counter$count = 84448;
	#10 counter$count = 84449;
	#10 counter$count = 84450;
	#10 counter$count = 84451;
	#10 counter$count = 84452;
	#10 counter$count = 84453;
	#10 counter$count = 84454;
	#10 counter$count = 84455;
	#10 counter$count = 84456;
	#10 counter$count = 84457;
	#10 counter$count = 84458;
	#10 counter$count = 84459;
	#10 counter$count = 84460;
	#10 counter$count = 84461;
	#10 counter$count = 84462;
	#10 counter$count = 84463;
	#10 counter$count = 84464;
	#10 counter$count = 84465;
	#10 counter$count = 84466;
	#10 counter$count = 84467;
	#10 counter$count = 84468;
	#10 counter$count = 84469;
	#10 counter$count = 84470;
	#10 counter$count = 84471;
	#10 counter$count = 84472;
	#10 counter$count = 84473;
	#10 counter$count = 84474;
	#10 counter$count = 84475;
	#10 counter$count = 84476;
	#10 counter$count = 84477;
	#10 counter$count = 84478;
	#10 counter$count = 84479;
	#10 counter$count = 84480;
	#10 counter$count = 84481;
	#10 counter$count = 84482;
	#10 counter$count = 84483;
	#10 counter$count = 84484;
	#10 counter$count = 84485;
	#10 counter$count = 84486;
	#10 counter$count = 84487;
	#10 counter$count = 84488;
	#10 counter$count = 84489;
	#10 counter$count = 84490;
	#10 counter$count = 84491;
	#10 counter$count = 84492;
	#10 counter$count = 84493;
	#10 counter$count = 84494;
	#10 counter$count = 84495;
	#10 counter$count = 84496;
	#10 counter$count = 84497;
	#10 counter$count = 84498;
	#10 counter$count = 84499;
	#10 counter$count = 84500;
	#10 counter$count = 84501;
	#10 counter$count = 84502;
	#10 counter$count = 84503;
	#10 counter$count = 84504;
	#10 counter$count = 84505;
	#10 counter$count = 84506;
	#10 counter$count = 84507;
	#10 counter$count = 84508;
	#10 counter$count = 84509;
	#10 counter$count = 84510;
	#10 counter$count = 84511;
	#10 counter$count = 84512;
	#10 counter$count = 84513;
	#10 counter$count = 84514;
	#10 counter$count = 84515;
	#10 counter$count = 84516;
	#10 counter$count = 84517;
	#10 counter$count = 84518;
	#10 counter$count = 84519;
	#10 counter$count = 84520;
	#10 counter$count = 84521;
	#10 counter$count = 84522;
	#10 counter$count = 84523;
	#10 counter$count = 84524;
	#10 counter$count = 84525;
	#10 counter$count = 84526;
	#10 counter$count = 84527;
	#10 counter$count = 84528;
	#10 counter$count = 84529;
	#10 counter$count = 84530;
	#10 counter$count = 84531;
	#10 counter$count = 84532;
	#10 counter$count = 84533;
	#10 counter$count = 84534;
	#10 counter$count = 84535;
	#10 counter$count = 84536;
	#10 counter$count = 84537;
	#10 counter$count = 84538;
	#10 counter$count = 84539;
	#10 counter$count = 84540;
	#10 counter$count = 84541;
	#10 counter$count = 84542;
	#10 counter$count = 84543;
	#10 counter$count = 84544;
	#10 counter$count = 84545;
	#10 counter$count = 84546;
	#10 counter$count = 84547;
	#10 counter$count = 84548;
	#10 counter$count = 84549;
	#10 counter$count = 84550;
	#10 counter$count = 84551;
	#10 counter$count = 84552;
	#10 counter$count = 84553;
	#10 counter$count = 84554;
	#10 counter$count = 84555;
	#10 counter$count = 84556;
	#10 counter$count = 84557;
	#10 counter$count = 84558;
	#10 counter$count = 84559;
	#10 counter$count = 84560;
	#10 counter$count = 84561;
	#10 counter$count = 84562;
	#10 counter$count = 84563;
	#10 counter$count = 84564;
	#10 counter$count = 84565;
	#10 counter$count = 84566;
	#10 counter$count = 84567;
	#10 counter$count = 84568;
	#10 counter$count = 84569;
	#10 counter$count = 84570;
	#10 counter$count = 84571;
	#10 counter$count = 84572;
	#10 counter$count = 84573;
	#10 counter$count = 84574;
	#10 counter$count = 84575;
	#10 counter$count = 84576;
	#10 counter$count = 84577;
	#10 counter$count = 84578;
	#10 counter$count = 84579;
	#10 counter$count = 84580;
	#10 counter$count = 84581;
	#10 counter$count = 84582;
	#10 counter$count = 84583;
	#10 counter$count = 84584;
	#10 counter$count = 84585;
	#10 counter$count = 84586;
	#10 counter$count = 84587;
	#10 counter$count = 84588;
	#10 counter$count = 84589;
	#10 counter$count = 84590;
	#10 counter$count = 84591;
	#10 counter$count = 84592;
	#10 counter$count = 84593;
	#10 counter$count = 84594;
	#10 counter$count = 84595;
	#10 counter$count = 84596;
	#10 counter$count = 84597;
	#10 counter$count = 84598;
	#10 counter$count = 84599;
	#10 counter$count = 84600;
	#10 counter$count = 84601;
	#10 counter$count = 84602;
	#10 counter$count = 84603;
	#10 counter$count = 84604;
	#10 counter$count = 84605;
	#10 counter$count = 84606;
	#10 counter$count = 84607;
	#10 counter$count = 84608;
	#10 counter$count = 84609;
	#10 counter$count = 84610;
	#10 counter$count = 84611;
	#10 counter$count = 84612;
	#10 counter$count = 84613;
	#10 counter$count = 84614;
	#10 counter$count = 84615;
	#10 counter$count = 84616;
	#10 counter$count = 84617;
	#10 counter$count = 84618;
	#10 counter$count = 84619;
	#10 counter$count = 84620;
	#10 counter$count = 84621;
	#10 counter$count = 84622;
	#10 counter$count = 84623;
	#10 counter$count = 84624;
	#10 counter$count = 84625;
	#10 counter$count = 84626;
	#10 counter$count = 84627;
	#10 counter$count = 84628;
	#10 counter$count = 84629;
	#10 counter$count = 84630;
	#10 counter$count = 84631;
	#10 counter$count = 84632;
	#10 counter$count = 84633;
	#10 counter$count = 84634;
	#10 counter$count = 84635;
	#10 counter$count = 84636;
	#10 counter$count = 84637;
	#10 counter$count = 84638;
	#10 counter$count = 84639;
	#10 counter$count = 84640;
	#10 counter$count = 84641;
	#10 counter$count = 84642;
	#10 counter$count = 84643;
	#10 counter$count = 84644;
	#10 counter$count = 84645;
	#10 counter$count = 84646;
	#10 counter$count = 84647;
	#10 counter$count = 84648;
	#10 counter$count = 84649;
	#10 counter$count = 84650;
	#10 counter$count = 84651;
	#10 counter$count = 84652;
	#10 counter$count = 84653;
	#10 counter$count = 84654;
	#10 counter$count = 84655;
	#10 counter$count = 84656;
	#10 counter$count = 84657;
	#10 counter$count = 84658;
	#10 counter$count = 84659;
	#10 counter$count = 84660;
	#10 counter$count = 84661;
	#10 counter$count = 84662;
	#10 counter$count = 84663;
	#10 counter$count = 84664;
	#10 counter$count = 84665;
	#10 counter$count = 84666;
	#10 counter$count = 84667;
	#10 counter$count = 84668;
	#10 counter$count = 84669;
	#10 counter$count = 84670;
	#10 counter$count = 84671;
	#10 counter$count = 84672;
	#10 counter$count = 84673;
	#10 counter$count = 84674;
	#10 counter$count = 84675;
	#10 counter$count = 84676;
	#10 counter$count = 84677;
	#10 counter$count = 84678;
	#10 counter$count = 84679;
	#10 counter$count = 84680;
	#10 counter$count = 84681;
	#10 counter$count = 84682;
	#10 counter$count = 84683;
	#10 counter$count = 84684;
	#10 counter$count = 84685;
	#10 counter$count = 84686;
	#10 counter$count = 84687;
	#10 counter$count = 84688;
	#10 counter$count = 84689;
	#10 counter$count = 84690;
	#10 counter$count = 84691;
	#10 counter$count = 84692;
	#10 counter$count = 84693;
	#10 counter$count = 84694;
	#10 counter$count = 84695;
	#10 counter$count = 84696;
	#10 counter$count = 84697;
	#10 counter$count = 84698;
	#10 counter$count = 84699;
	#10 counter$count = 84700;
	#10 counter$count = 84701;
	#10 counter$count = 84702;
	#10 counter$count = 84703;
	#10 counter$count = 84704;
	#10 counter$count = 84705;
	#10 counter$count = 84706;
	#10 counter$count = 84707;
	#10 counter$count = 84708;
	#10 counter$count = 84709;
	#10 counter$count = 84710;
	#10 counter$count = 84711;
	#10 counter$count = 84712;
	#10 counter$count = 84713;
	#10 counter$count = 84714;
	#10 counter$count = 84715;
	#10 counter$count = 84716;
	#10 counter$count = 84717;
	#10 counter$count = 84718;
	#10 counter$count = 84719;
	#10 counter$count = 84720;
	#10 counter$count = 84721;
	#10 counter$count = 84722;
	#10 counter$count = 84723;
	#10 counter$count = 84724;
	#10 counter$count = 84725;
	#10 counter$count = 84726;
	#10 counter$count = 84727;
	#10 counter$count = 84728;
	#10 counter$count = 84729;
	#10 counter$count = 84730;
	#10 counter$count = 84731;
	#10 counter$count = 84732;
	#10 counter$count = 84733;
	#10 counter$count = 84734;
	#10 counter$count = 84735;
	#10 counter$count = 84736;
	#10 counter$count = 84737;
	#10 counter$count = 84738;
	#10 counter$count = 84739;
	#10 counter$count = 84740;
	#10 counter$count = 84741;
	#10 counter$count = 84742;
	#10 counter$count = 84743;
	#10 counter$count = 84744;
	#10 counter$count = 84745;
	#10 counter$count = 84746;
	#10 counter$count = 84747;
	#10 counter$count = 84748;
	#10 counter$count = 84749;
	#10 counter$count = 84750;
	#10 counter$count = 84751;
	#10 counter$count = 84752;
	#10 counter$count = 84753;
	#10 counter$count = 84754;
	#10 counter$count = 84755;
	#10 counter$count = 84756;
	#10 counter$count = 84757;
	#10 counter$count = 84758;
	#10 counter$count = 84759;
	#10 counter$count = 84760;
	#10 counter$count = 84761;
	#10 counter$count = 84762;
	#10 counter$count = 84763;
	#10 counter$count = 84764;
	#10 counter$count = 84765;
	#10 counter$count = 84766;
	#10 counter$count = 84767;
	#10 counter$count = 84768;
	#10 counter$count = 84769;
	#10 counter$count = 84770;
	#10 counter$count = 84771;
	#10 counter$count = 84772;
	#10 counter$count = 84773;
	#10 counter$count = 84774;
	#10 counter$count = 84775;
	#10 counter$count = 84776;
	#10 counter$count = 84777;
	#10 counter$count = 84778;
	#10 counter$count = 84779;
	#10 counter$count = 84780;
	#10 counter$count = 84781;
	#10 counter$count = 84782;
	#10 counter$count = 84783;
	#10 counter$count = 84784;
	#10 counter$count = 84785;
	#10 counter$count = 84786;
	#10 counter$count = 84787;
	#10 counter$count = 84788;
	#10 counter$count = 84789;
	#10 counter$count = 84790;
	#10 counter$count = 84791;
	#10 counter$count = 84792;
	#10 counter$count = 84793;
	#10 counter$count = 84794;
	#10 counter$count = 84795;
	#10 counter$count = 84796;
	#10 counter$count = 84797;
	#10 counter$count = 84798;
	#10 counter$count = 84799;
	#10 counter$count = 84800;
	#10 counter$count = 84801;
	#10 counter$count = 84802;
	#10 counter$count = 84803;
	#10 counter$count = 84804;
	#10 counter$count = 84805;
	#10 counter$count = 84806;
	#10 counter$count = 84807;
	#10 counter$count = 84808;
	#10 counter$count = 84809;
	#10 counter$count = 84810;
	#10 counter$count = 84811;
	#10 counter$count = 84812;
	#10 counter$count = 84813;
	#10 counter$count = 84814;
	#10 counter$count = 84815;
	#10 counter$count = 84816;
	#10 counter$count = 84817;
	#10 counter$count = 84818;
	#10 counter$count = 84819;
	#10 counter$count = 84820;
	#10 counter$count = 84821;
	#10 counter$count = 84822;
	#10 counter$count = 84823;
	#10 counter$count = 84824;
	#10 counter$count = 84825;
	#10 counter$count = 84826;
	#10 counter$count = 84827;
	#10 counter$count = 84828;
	#10 counter$count = 84829;
	#10 counter$count = 84830;
	#10 counter$count = 84831;
	#10 counter$count = 84832;
	#10 counter$count = 84833;
	#10 counter$count = 84834;
	#10 counter$count = 84835;
	#10 counter$count = 84836;
	#10 counter$count = 84837;
	#10 counter$count = 84838;
	#10 counter$count = 84839;
	#10 counter$count = 84840;
	#10 counter$count = 84841;
	#10 counter$count = 84842;
	#10 counter$count = 84843;
	#10 counter$count = 84844;
	#10 counter$count = 84845;
	#10 counter$count = 84846;
	#10 counter$count = 84847;
	#10 counter$count = 84848;
	#10 counter$count = 84849;
	#10 counter$count = 84850;
	#10 counter$count = 84851;
	#10 counter$count = 84852;
	#10 counter$count = 84853;
	#10 counter$count = 84854;
	#10 counter$count = 84855;
	#10 counter$count = 84856;
	#10 counter$count = 84857;
	#10 counter$count = 84858;
	#10 counter$count = 84859;
	#10 counter$count = 84860;
	#10 counter$count = 84861;
	#10 counter$count = 84862;
	#10 counter$count = 84863;
	#10 counter$count = 84864;
	#10 counter$count = 84865;
	#10 counter$count = 84866;
	#10 counter$count = 84867;
	#10 counter$count = 84868;
	#10 counter$count = 84869;
	#10 counter$count = 84870;
	#10 counter$count = 84871;
	#10 counter$count = 84872;
	#10 counter$count = 84873;
	#10 counter$count = 84874;
	#10 counter$count = 84875;
	#10 counter$count = 84876;
	#10 counter$count = 84877;
	#10 counter$count = 84878;
	#10 counter$count = 84879;
	#10 counter$count = 84880;
	#10 counter$count = 84881;
	#10 counter$count = 84882;
	#10 counter$count = 84883;
	#10 counter$count = 84884;
	#10 counter$count = 84885;
	#10 counter$count = 84886;
	#10 counter$count = 84887;
	#10 counter$count = 84888;
	#10 counter$count = 84889;
	#10 counter$count = 84890;
	#10 counter$count = 84891;
	#10 counter$count = 84892;
	#10 counter$count = 84893;
	#10 counter$count = 84894;
	#10 counter$count = 84895;
	#10 counter$count = 84896;
	#10 counter$count = 84897;
	#10 counter$count = 84898;
	#10 counter$count = 84899;
	#10 counter$count = 84900;
	#10 counter$count = 84901;
	#10 counter$count = 84902;
	#10 counter$count = 84903;
	#10 counter$count = 84904;
	#10 counter$count = 84905;
	#10 counter$count = 84906;
	#10 counter$count = 84907;
	#10 counter$count = 84908;
	#10 counter$count = 84909;
	#10 counter$count = 84910;
	#10 counter$count = 84911;
	#10 counter$count = 84912;
	#10 counter$count = 84913;
	#10 counter$count = 84914;
	#10 counter$count = 84915;
	#10 counter$count = 84916;
	#10 counter$count = 84917;
	#10 counter$count = 84918;
	#10 counter$count = 84919;
	#10 counter$count = 84920;
	#10 counter$count = 84921;
	#10 counter$count = 84922;
	#10 counter$count = 84923;
	#10 counter$count = 84924;
	#10 counter$count = 84925;
	#10 counter$count = 84926;
	#10 counter$count = 84927;
	#10 counter$count = 84928;
	#10 counter$count = 84929;
	#10 counter$count = 84930;
	#10 counter$count = 84931;
	#10 counter$count = 84932;
	#10 counter$count = 84933;
	#10 counter$count = 84934;
	#10 counter$count = 84935;
	#10 counter$count = 84936;
	#10 counter$count = 84937;
	#10 counter$count = 84938;
	#10 counter$count = 84939;
	#10 counter$count = 84940;
	#10 counter$count = 84941;
	#10 counter$count = 84942;
	#10 counter$count = 84943;
	#10 counter$count = 84944;
	#10 counter$count = 84945;
	#10 counter$count = 84946;
	#10 counter$count = 84947;
	#10 counter$count = 84948;
	#10 counter$count = 84949;
	#10 counter$count = 84950;
	#10 counter$count = 84951;
	#10 counter$count = 84952;
	#10 counter$count = 84953;
	#10 counter$count = 84954;
	#10 counter$count = 84955;
	#10 counter$count = 84956;
	#10 counter$count = 84957;
	#10 counter$count = 84958;
	#10 counter$count = 84959;
	#10 counter$count = 84960;
	#10 counter$count = 84961;
	#10 counter$count = 84962;
	#10 counter$count = 84963;
	#10 counter$count = 84964;
	#10 counter$count = 84965;
	#10 counter$count = 84966;
	#10 counter$count = 84967;
	#10 counter$count = 84968;
	#10 counter$count = 84969;
	#10 counter$count = 84970;
	#10 counter$count = 84971;
	#10 counter$count = 84972;
	#10 counter$count = 84973;
	#10 counter$count = 84974;
	#10 counter$count = 84975;
	#10 counter$count = 84976;
	#10 counter$count = 84977;
	#10 counter$count = 84978;
	#10 counter$count = 84979;
	#10 counter$count = 84980;
	#10 counter$count = 84981;
	#10 counter$count = 84982;
	#10 counter$count = 84983;
	#10 counter$count = 84984;
	#10 counter$count = 84985;
	#10 counter$count = 84986;
	#10 counter$count = 84987;
	#10 counter$count = 84988;
	#10 counter$count = 84989;
	#10 counter$count = 84990;
	#10 counter$count = 84991;
	#10 counter$count = 84992;
	#10 counter$count = 84993;
	#10 counter$count = 84994;
	#10 counter$count = 84995;
	#10 counter$count = 84996;
	#10 counter$count = 84997;
	#10 counter$count = 84998;
	#10 counter$count = 84999;
	#10 counter$count = 85000;
	#10 counter$count = 85001;
	#10 counter$count = 85002;
	#10 counter$count = 85003;
	#10 counter$count = 85004;
	#10 counter$count = 85005;
	#10 counter$count = 85006;
	#10 counter$count = 85007;
	#10 counter$count = 85008;
	#10 counter$count = 85009;
	#10 counter$count = 85010;
	#10 counter$count = 85011;
	#10 counter$count = 85012;
	#10 counter$count = 85013;
	#10 counter$count = 85014;
	#10 counter$count = 85015;
	#10 counter$count = 85016;
	#10 counter$count = 85017;
	#10 counter$count = 85018;
	#10 counter$count = 85019;
	#10 counter$count = 85020;
	#10 counter$count = 85021;
	#10 counter$count = 85022;
	#10 counter$count = 85023;
	#10 counter$count = 85024;
	#10 counter$count = 85025;
	#10 counter$count = 85026;
	#10 counter$count = 85027;
	#10 counter$count = 85028;
	#10 counter$count = 85029;
	#10 counter$count = 85030;
	#10 counter$count = 85031;
	#10 counter$count = 85032;
	#10 counter$count = 85033;
	#10 counter$count = 85034;
	#10 counter$count = 85035;
	#10 counter$count = 85036;
	#10 counter$count = 85037;
	#10 counter$count = 85038;
	#10 counter$count = 85039;
	#10 counter$count = 85040;
	#10 counter$count = 85041;
	#10 counter$count = 85042;
	#10 counter$count = 85043;
	#10 counter$count = 85044;
	#10 counter$count = 85045;
	#10 counter$count = 85046;
	#10 counter$count = 85047;
	#10 counter$count = 85048;
	#10 counter$count = 85049;
	#10 counter$count = 85050;
	#10 counter$count = 85051;
	#10 counter$count = 85052;
	#10 counter$count = 85053;
	#10 counter$count = 85054;
	#10 counter$count = 85055;
	#10 counter$count = 85056;
	#10 counter$count = 85057;
	#10 counter$count = 85058;
	#10 counter$count = 85059;
	#10 counter$count = 85060;
	#10 counter$count = 85061;
	#10 counter$count = 85062;
	#10 counter$count = 85063;
	#10 counter$count = 85064;
	#10 counter$count = 85065;
	#10 counter$count = 85066;
	#10 counter$count = 85067;
	#10 counter$count = 85068;
	#10 counter$count = 85069;
	#10 counter$count = 85070;
	#10 counter$count = 85071;
	#10 counter$count = 85072;
	#10 counter$count = 85073;
	#10 counter$count = 85074;
	#10 counter$count = 85075;
	#10 counter$count = 85076;
	#10 counter$count = 85077;
	#10 counter$count = 85078;
	#10 counter$count = 85079;
	#10 counter$count = 85080;
	#10 counter$count = 85081;
	#10 counter$count = 85082;
	#10 counter$count = 85083;
	#10 counter$count = 85084;
	#10 counter$count = 85085;
	#10 counter$count = 85086;
	#10 counter$count = 85087;
	#10 counter$count = 85088;
	#10 counter$count = 85089;
	#10 counter$count = 85090;
	#10 counter$count = 85091;
	#10 counter$count = 85092;
	#10 counter$count = 85093;
	#10 counter$count = 85094;
	#10 counter$count = 85095;
	#10 counter$count = 85096;
	#10 counter$count = 85097;
	#10 counter$count = 85098;
	#10 counter$count = 85099;
	#10 counter$count = 85100;
	#10 counter$count = 85101;
	#10 counter$count = 85102;
	#10 counter$count = 85103;
	#10 counter$count = 85104;
	#10 counter$count = 85105;
	#10 counter$count = 85106;
	#10 counter$count = 85107;
	#10 counter$count = 85108;
	#10 counter$count = 85109;
	#10 counter$count = 85110;
	#10 counter$count = 85111;
	#10 counter$count = 85112;
	#10 counter$count = 85113;
	#10 counter$count = 85114;
	#10 counter$count = 85115;
	#10 counter$count = 85116;
	#10 counter$count = 85117;
	#10 counter$count = 85118;
	#10 counter$count = 85119;
	#10 counter$count = 85120;
	#10 counter$count = 85121;
	#10 counter$count = 85122;
	#10 counter$count = 85123;
	#10 counter$count = 85124;
	#10 counter$count = 85125;
	#10 counter$count = 85126;
	#10 counter$count = 85127;
	#10 counter$count = 85128;
	#10 counter$count = 85129;
	#10 counter$count = 85130;
	#10 counter$count = 85131;
	#10 counter$count = 85132;
	#10 counter$count = 85133;
	#10 counter$count = 85134;
	#10 counter$count = 85135;
	#10 counter$count = 85136;
	#10 counter$count = 85137;
	#10 counter$count = 85138;
	#10 counter$count = 85139;
	#10 counter$count = 85140;
	#10 counter$count = 85141;
	#10 counter$count = 85142;
	#10 counter$count = 85143;
	#10 counter$count = 85144;
	#10 counter$count = 85145;
	#10 counter$count = 85146;
	#10 counter$count = 85147;
	#10 counter$count = 85148;
	#10 counter$count = 85149;
	#10 counter$count = 85150;
	#10 counter$count = 85151;
	#10 counter$count = 85152;
	#10 counter$count = 85153;
	#10 counter$count = 85154;
	#10 counter$count = 85155;
	#10 counter$count = 85156;
	#10 counter$count = 85157;
	#10 counter$count = 85158;
	#10 counter$count = 85159;
	#10 counter$count = 85160;
	#10 counter$count = 85161;
	#10 counter$count = 85162;
	#10 counter$count = 85163;
	#10 counter$count = 85164;
	#10 counter$count = 85165;
	#10 counter$count = 85166;
	#10 counter$count = 85167;
	#10 counter$count = 85168;
	#10 counter$count = 85169;
	#10 counter$count = 85170;
	#10 counter$count = 85171;
	#10 counter$count = 85172;
	#10 counter$count = 85173;
	#10 counter$count = 85174;
	#10 counter$count = 85175;
	#10 counter$count = 85176;
	#10 counter$count = 85177;
	#10 counter$count = 85178;
	#10 counter$count = 85179;
	#10 counter$count = 85180;
	#10 counter$count = 85181;
	#10 counter$count = 85182;
	#10 counter$count = 85183;
	#10 counter$count = 85184;
	#10 counter$count = 85185;
	#10 counter$count = 85186;
	#10 counter$count = 85187;
	#10 counter$count = 85188;
	#10 counter$count = 85189;
	#10 counter$count = 85190;
	#10 counter$count = 85191;
	#10 counter$count = 85192;
	#10 counter$count = 85193;
	#10 counter$count = 85194;
	#10 counter$count = 85195;
	#10 counter$count = 85196;
	#10 counter$count = 85197;
	#10 counter$count = 85198;
	#10 counter$count = 85199;
	#10 counter$count = 85200;
	#10 counter$count = 85201;
	#10 counter$count = 85202;
	#10 counter$count = 85203;
	#10 counter$count = 85204;
	#10 counter$count = 85205;
	#10 counter$count = 85206;
	#10 counter$count = 85207;
	#10 counter$count = 85208;
	#10 counter$count = 85209;
	#10 counter$count = 85210;
	#10 counter$count = 85211;
	#10 counter$count = 85212;
	#10 counter$count = 85213;
	#10 counter$count = 85214;
	#10 counter$count = 85215;
	#10 counter$count = 85216;
	#10 counter$count = 85217;
	#10 counter$count = 85218;
	#10 counter$count = 85219;
	#10 counter$count = 85220;
	#10 counter$count = 85221;
	#10 counter$count = 85222;
	#10 counter$count = 85223;
	#10 counter$count = 85224;
	#10 counter$count = 85225;
	#10 counter$count = 85226;
	#10 counter$count = 85227;
	#10 counter$count = 85228;
	#10 counter$count = 85229;
	#10 counter$count = 85230;
	#10 counter$count = 85231;
	#10 counter$count = 85232;
	#10 counter$count = 85233;
	#10 counter$count = 85234;
	#10 counter$count = 85235;
	#10 counter$count = 85236;
	#10 counter$count = 85237;
	#10 counter$count = 85238;
	#10 counter$count = 85239;
	#10 counter$count = 85240;
	#10 counter$count = 85241;
	#10 counter$count = 85242;
	#10 counter$count = 85243;
	#10 counter$count = 85244;
	#10 counter$count = 85245;
	#10 counter$count = 85246;
	#10 counter$count = 85247;
	#10 counter$count = 85248;
	#10 counter$count = 85249;
	#10 counter$count = 85250;
	#10 counter$count = 85251;
	#10 counter$count = 85252;
	#10 counter$count = 85253;
	#10 counter$count = 85254;
	#10 counter$count = 85255;
	#10 counter$count = 85256;
	#10 counter$count = 85257;
	#10 counter$count = 85258;
	#10 counter$count = 85259;
	#10 counter$count = 85260;
	#10 counter$count = 85261;
	#10 counter$count = 85262;
	#10 counter$count = 85263;
	#10 counter$count = 85264;
	#10 counter$count = 85265;
	#10 counter$count = 85266;
	#10 counter$count = 85267;
	#10 counter$count = 85268;
	#10 counter$count = 85269;
	#10 counter$count = 85270;
	#10 counter$count = 85271;
	#10 counter$count = 85272;
	#10 counter$count = 85273;
	#10 counter$count = 85274;
	#10 counter$count = 85275;
	#10 counter$count = 85276;
	#10 counter$count = 85277;
	#10 counter$count = 85278;
	#10 counter$count = 85279;
	#10 counter$count = 85280;
	#10 counter$count = 85281;
	#10 counter$count = 85282;
	#10 counter$count = 85283;
	#10 counter$count = 85284;
	#10 counter$count = 85285;
	#10 counter$count = 85286;
	#10 counter$count = 85287;
	#10 counter$count = 85288;
	#10 counter$count = 85289;
	#10 counter$count = 85290;
	#10 counter$count = 85291;
	#10 counter$count = 85292;
	#10 counter$count = 85293;
	#10 counter$count = 85294;
	#10 counter$count = 85295;
	#10 counter$count = 85296;
	#10 counter$count = 85297;
	#10 counter$count = 85298;
	#10 counter$count = 85299;
	#10 counter$count = 85300;
	#10 counter$count = 85301;
	#10 counter$count = 85302;
	#10 counter$count = 85303;
	#10 counter$count = 85304;
	#10 counter$count = 85305;
	#10 counter$count = 85306;
	#10 counter$count = 85307;
	#10 counter$count = 85308;
	#10 counter$count = 85309;
	#10 counter$count = 85310;
	#10 counter$count = 85311;
	#10 counter$count = 85312;
	#10 counter$count = 85313;
	#10 counter$count = 85314;
	#10 counter$count = 85315;
	#10 counter$count = 85316;
	#10 counter$count = 85317;
	#10 counter$count = 85318;
	#10 counter$count = 85319;
	#10 counter$count = 85320;
	#10 counter$count = 85321;
	#10 counter$count = 85322;
	#10 counter$count = 85323;
	#10 counter$count = 85324;
	#10 counter$count = 85325;
	#10 counter$count = 85326;
	#10 counter$count = 85327;
	#10 counter$count = 85328;
	#10 counter$count = 85329;
	#10 counter$count = 85330;
	#10 counter$count = 85331;
	#10 counter$count = 85332;
	#10 counter$count = 85333;
	#10 counter$count = 85334;
	#10 counter$count = 85335;
	#10 counter$count = 85336;
	#10 counter$count = 85337;
	#10 counter$count = 85338;
	#10 counter$count = 85339;
	#10 counter$count = 85340;
	#10 counter$count = 85341;
	#10 counter$count = 85342;
	#10 counter$count = 85343;
	#10 counter$count = 85344;
	#10 counter$count = 85345;
	#10 counter$count = 85346;
	#10 counter$count = 85347;
	#10 counter$count = 85348;
	#10 counter$count = 85349;
	#10 counter$count = 85350;
	#10 counter$count = 85351;
	#10 counter$count = 85352;
	#10 counter$count = 85353;
	#10 counter$count = 85354;
	#10 counter$count = 85355;
	#10 counter$count = 85356;
	#10 counter$count = 85357;
	#10 counter$count = 85358;
	#10 counter$count = 85359;
	#10 counter$count = 85360;
	#10 counter$count = 85361;
	#10 counter$count = 85362;
	#10 counter$count = 85363;
	#10 counter$count = 85364;
	#10 counter$count = 85365;
	#10 counter$count = 85366;
	#10 counter$count = 85367;
	#10 counter$count = 85368;
	#10 counter$count = 85369;
	#10 counter$count = 85370;
	#10 counter$count = 85371;
	#10 counter$count = 85372;
	#10 counter$count = 85373;
	#10 counter$count = 85374;
	#10 counter$count = 85375;
	#10 counter$count = 85376;
	#10 counter$count = 85377;
	#10 counter$count = 85378;
	#10 counter$count = 85379;
	#10 counter$count = 85380;
	#10 counter$count = 85381;
	#10 counter$count = 85382;
	#10 counter$count = 85383;
	#10 counter$count = 85384;
	#10 counter$count = 85385;
	#10 counter$count = 85386;
	#10 counter$count = 85387;
	#10 counter$count = 85388;
	#10 counter$count = 85389;
	#10 counter$count = 85390;
	#10 counter$count = 85391;
	#10 counter$count = 85392;
	#10 counter$count = 85393;
	#10 counter$count = 85394;
	#10 counter$count = 85395;
	#10 counter$count = 85396;
	#10 counter$count = 85397;
	#10 counter$count = 85398;
	#10 counter$count = 85399;
	#10 counter$count = 85400;
	#10 counter$count = 85401;
	#10 counter$count = 85402;
	#10 counter$count = 85403;
	#10 counter$count = 85404;
	#10 counter$count = 85405;
	#10 counter$count = 85406;
	#10 counter$count = 85407;
	#10 counter$count = 85408;
	#10 counter$count = 85409;
	#10 counter$count = 85410;
	#10 counter$count = 85411;
	#10 counter$count = 85412;
	#10 counter$count = 85413;
	#10 counter$count = 85414;
	#10 counter$count = 85415;
	#10 counter$count = 85416;
	#10 counter$count = 85417;
	#10 counter$count = 85418;
	#10 counter$count = 85419;
	#10 counter$count = 85420;
	#10 counter$count = 85421;
	#10 counter$count = 85422;
	#10 counter$count = 85423;
	#10 counter$count = 85424;
	#10 counter$count = 85425;
	#10 counter$count = 85426;
	#10 counter$count = 85427;
	#10 counter$count = 85428;
	#10 counter$count = 85429;
	#10 counter$count = 85430;
	#10 counter$count = 85431;
	#10 counter$count = 85432;
	#10 counter$count = 85433;
	#10 counter$count = 85434;
	#10 counter$count = 85435;
	#10 counter$count = 85436;
	#10 counter$count = 85437;
	#10 counter$count = 85438;
	#10 counter$count = 85439;
	#10 counter$count = 85440;
	#10 counter$count = 85441;
	#10 counter$count = 85442;
	#10 counter$count = 85443;
	#10 counter$count = 85444;
	#10 counter$count = 85445;
	#10 counter$count = 85446;
	#10 counter$count = 85447;
	#10 counter$count = 85448;
	#10 counter$count = 85449;
	#10 counter$count = 85450;
	#10 counter$count = 85451;
	#10 counter$count = 85452;
	#10 counter$count = 85453;
	#10 counter$count = 85454;
	#10 counter$count = 85455;
	#10 counter$count = 85456;
	#10 counter$count = 85457;
	#10 counter$count = 85458;
	#10 counter$count = 85459;
	#10 counter$count = 85460;
	#10 counter$count = 85461;
	#10 counter$count = 85462;
	#10 counter$count = 85463;
	#10 counter$count = 85464;
	#10 counter$count = 85465;
	#10 counter$count = 85466;
	#10 counter$count = 85467;
	#10 counter$count = 85468;
	#10 counter$count = 85469;
	#10 counter$count = 85470;
	#10 counter$count = 85471;
	#10 counter$count = 85472;
	#10 counter$count = 85473;
	#10 counter$count = 85474;
	#10 counter$count = 85475;
	#10 counter$count = 85476;
	#10 counter$count = 85477;
	#10 counter$count = 85478;
	#10 counter$count = 85479;
	#10 counter$count = 85480;
	#10 counter$count = 85481;
	#10 counter$count = 85482;
	#10 counter$count = 85483;
	#10 counter$count = 85484;
	#10 counter$count = 85485;
	#10 counter$count = 85486;
	#10 counter$count = 85487;
	#10 counter$count = 85488;
	#10 counter$count = 85489;
	#10 counter$count = 85490;
	#10 counter$count = 85491;
	#10 counter$count = 85492;
	#10 counter$count = 85493;
	#10 counter$count = 85494;
	#10 counter$count = 85495;
	#10 counter$count = 85496;
	#10 counter$count = 85497;
	#10 counter$count = 85498;
	#10 counter$count = 85499;
	#10 counter$count = 85500;
	#10 counter$count = 85501;
	#10 counter$count = 85502;
	#10 counter$count = 85503;
	#10 counter$count = 85504;
	#10 counter$count = 85505;
	#10 counter$count = 85506;
	#10 counter$count = 85507;
	#10 counter$count = 85508;
	#10 counter$count = 85509;
	#10 counter$count = 85510;
	#10 counter$count = 85511;
	#10 counter$count = 85512;
	#10 counter$count = 85513;
	#10 counter$count = 85514;
	#10 counter$count = 85515;
	#10 counter$count = 85516;
	#10 counter$count = 85517;
	#10 counter$count = 85518;
	#10 counter$count = 85519;
	#10 counter$count = 85520;
	#10 counter$count = 85521;
	#10 counter$count = 85522;
	#10 counter$count = 85523;
	#10 counter$count = 85524;
	#10 counter$count = 85525;
	#10 counter$count = 85526;
	#10 counter$count = 85527;
	#10 counter$count = 85528;
	#10 counter$count = 85529;
	#10 counter$count = 85530;
	#10 counter$count = 85531;
	#10 counter$count = 85532;
	#10 counter$count = 85533;
	#10 counter$count = 85534;
	#10 counter$count = 85535;
	#10 counter$count = 85536;
	#10 counter$count = 85537;
	#10 counter$count = 85538;
	#10 counter$count = 85539;
	#10 counter$count = 85540;
	#10 counter$count = 85541;
	#10 counter$count = 85542;
	#10 counter$count = 85543;
	#10 counter$count = 85544;
	#10 counter$count = 85545;
	#10 counter$count = 85546;
	#10 counter$count = 85547;
	#10 counter$count = 85548;
	#10 counter$count = 85549;
	#10 counter$count = 85550;
	#10 counter$count = 85551;
	#10 counter$count = 85552;
	#10 counter$count = 85553;
	#10 counter$count = 85554;
	#10 counter$count = 85555;
	#10 counter$count = 85556;
	#10 counter$count = 85557;
	#10 counter$count = 85558;
	#10 counter$count = 85559;
	#10 counter$count = 85560;
	#10 counter$count = 85561;
	#10 counter$count = 85562;
	#10 counter$count = 85563;
	#10 counter$count = 85564;
	#10 counter$count = 85565;
	#10 counter$count = 85566;
	#10 counter$count = 85567;
	#10 counter$count = 85568;
	#10 counter$count = 85569;
	#10 counter$count = 85570;
	#10 counter$count = 85571;
	#10 counter$count = 85572;
	#10 counter$count = 85573;
	#10 counter$count = 85574;
	#10 counter$count = 85575;
	#10 counter$count = 85576;
	#10 counter$count = 85577;
	#10 counter$count = 85578;
	#10 counter$count = 85579;
	#10 counter$count = 85580;
	#10 counter$count = 85581;
	#10 counter$count = 85582;
	#10 counter$count = 85583;
	#10 counter$count = 85584;
	#10 counter$count = 85585;
	#10 counter$count = 85586;
	#10 counter$count = 85587;
	#10 counter$count = 85588;
	#10 counter$count = 85589;
	#10 counter$count = 85590;
	#10 counter$count = 85591;
	#10 counter$count = 85592;
	#10 counter$count = 85593;
	#10 counter$count = 85594;
	#10 counter$count = 85595;
	#10 counter$count = 85596;
	#10 counter$count = 85597;
	#10 counter$count = 85598;
	#10 counter$count = 85599;
	#10 counter$count = 85600;
	#10 counter$count = 85601;
	#10 counter$count = 85602;
	#10 counter$count = 85603;
	#10 counter$count = 85604;
	#10 counter$count = 85605;
	#10 counter$count = 85606;
	#10 counter$count = 85607;
	#10 counter$count = 85608;
	#10 counter$count = 85609;
	#10 counter$count = 85610;
	#10 counter$count = 85611;
	#10 counter$count = 85612;
	#10 counter$count = 85613;
	#10 counter$count = 85614;
	#10 counter$count = 85615;
	#10 counter$count = 85616;
	#10 counter$count = 85617;
	#10 counter$count = 85618;
	#10 counter$count = 85619;
	#10 counter$count = 85620;
	#10 counter$count = 85621;
	#10 counter$count = 85622;
	#10 counter$count = 85623;
	#10 counter$count = 85624;
	#10 counter$count = 85625;
	#10 counter$count = 85626;
	#10 counter$count = 85627;
	#10 counter$count = 85628;
	#10 counter$count = 85629;
	#10 counter$count = 85630;
	#10 counter$count = 85631;
	#10 counter$count = 85632;
	#10 counter$count = 85633;
	#10 counter$count = 85634;
	#10 counter$count = 85635;
	#10 counter$count = 85636;
	#10 counter$count = 85637;
	#10 counter$count = 85638;
	#10 counter$count = 85639;
	#10 counter$count = 85640;
	#10 counter$count = 85641;
	#10 counter$count = 85642;
	#10 counter$count = 85643;
	#10 counter$count = 85644;
	#10 counter$count = 85645;
	#10 counter$count = 85646;
	#10 counter$count = 85647;
	#10 counter$count = 85648;
	#10 counter$count = 85649;
	#10 counter$count = 85650;
	#10 counter$count = 85651;
	#10 counter$count = 85652;
	#10 counter$count = 85653;
	#10 counter$count = 85654;
	#10 counter$count = 85655;
	#10 counter$count = 85656;
	#10 counter$count = 85657;
	#10 counter$count = 85658;
	#10 counter$count = 85659;
	#10 counter$count = 85660;
	#10 counter$count = 85661;
	#10 counter$count = 85662;
	#10 counter$count = 85663;
	#10 counter$count = 85664;
	#10 counter$count = 85665;
	#10 counter$count = 85666;
	#10 counter$count = 85667;
	#10 counter$count = 85668;
	#10 counter$count = 85669;
	#10 counter$count = 85670;
	#10 counter$count = 85671;
	#10 counter$count = 85672;
	#10 counter$count = 85673;
	#10 counter$count = 85674;
	#10 counter$count = 85675;
	#10 counter$count = 85676;
	#10 counter$count = 85677;
	#10 counter$count = 85678;
	#10 counter$count = 85679;
	#10 counter$count = 85680;
	#10 counter$count = 85681;
	#10 counter$count = 85682;
	#10 counter$count = 85683;
	#10 counter$count = 85684;
	#10 counter$count = 85685;
	#10 counter$count = 85686;
	#10 counter$count = 85687;
	#10 counter$count = 85688;
	#10 counter$count = 85689;
	#10 counter$count = 85690;
	#10 counter$count = 85691;
	#10 counter$count = 85692;
	#10 counter$count = 85693;
	#10 counter$count = 85694;
	#10 counter$count = 85695;
	#10 counter$count = 85696;
	#10 counter$count = 85697;
	#10 counter$count = 85698;
	#10 counter$count = 85699;
	#10 counter$count = 85700;
	#10 counter$count = 85701;
	#10 counter$count = 85702;
	#10 counter$count = 85703;
	#10 counter$count = 85704;
	#10 counter$count = 85705;
	#10 counter$count = 85706;
	#10 counter$count = 85707;
	#10 counter$count = 85708;
	#10 counter$count = 85709;
	#10 counter$count = 85710;
	#10 counter$count = 85711;
	#10 counter$count = 85712;
	#10 counter$count = 85713;
	#10 counter$count = 85714;
	#10 counter$count = 85715;
	#10 counter$count = 85716;
	#10 counter$count = 85717;
	#10 counter$count = 85718;
	#10 counter$count = 85719;
	#10 counter$count = 85720;
	#10 counter$count = 85721;
	#10 counter$count = 85722;
	#10 counter$count = 85723;
	#10 counter$count = 85724;
	#10 counter$count = 85725;
	#10 counter$count = 85726;
	#10 counter$count = 85727;
	#10 counter$count = 85728;
	#10 counter$count = 85729;
	#10 counter$count = 85730;
	#10 counter$count = 85731;
	#10 counter$count = 85732;
	#10 counter$count = 85733;
	#10 counter$count = 85734;
	#10 counter$count = 85735;
	#10 counter$count = 85736;
	#10 counter$count = 85737;
	#10 counter$count = 85738;
	#10 counter$count = 85739;
	#10 counter$count = 85740;
	#10 counter$count = 85741;
	#10 counter$count = 85742;
	#10 counter$count = 85743;
	#10 counter$count = 85744;
	#10 counter$count = 85745;
	#10 counter$count = 85746;
	#10 counter$count = 85747;
	#10 counter$count = 85748;
	#10 counter$count = 85749;
	#10 counter$count = 85750;
	#10 counter$count = 85751;
	#10 counter$count = 85752;
	#10 counter$count = 85753;
	#10 counter$count = 85754;
	#10 counter$count = 85755;
	#10 counter$count = 85756;
	#10 counter$count = 85757;
	#10 counter$count = 85758;
	#10 counter$count = 85759;
	#10 counter$count = 85760;
	#10 counter$count = 85761;
	#10 counter$count = 85762;
	#10 counter$count = 85763;
	#10 counter$count = 85764;
	#10 counter$count = 85765;
	#10 counter$count = 85766;
	#10 counter$count = 85767;
	#10 counter$count = 85768;
	#10 counter$count = 85769;
	#10 counter$count = 85770;
	#10 counter$count = 85771;
	#10 counter$count = 85772;
	#10 counter$count = 85773;
	#10 counter$count = 85774;
	#10 counter$count = 85775;
	#10 counter$count = 85776;
	#10 counter$count = 85777;
	#10 counter$count = 85778;
	#10 counter$count = 85779;
	#10 counter$count = 85780;
	#10 counter$count = 85781;
	#10 counter$count = 85782;
	#10 counter$count = 85783;
	#10 counter$count = 85784;
	#10 counter$count = 85785;
	#10 counter$count = 85786;
	#10 counter$count = 85787;
	#10 counter$count = 85788;
	#10 counter$count = 85789;
	#10 counter$count = 85790;
	#10 counter$count = 85791;
	#10 counter$count = 85792;
	#10 counter$count = 85793;
	#10 counter$count = 85794;
	#10 counter$count = 85795;
	#10 counter$count = 85796;
	#10 counter$count = 85797;
	#10 counter$count = 85798;
	#10 counter$count = 85799;
	#10 counter$count = 85800;
	#10 counter$count = 85801;
	#10 counter$count = 85802;
	#10 counter$count = 85803;
	#10 counter$count = 85804;
	#10 counter$count = 85805;
	#10 counter$count = 85806;
	#10 counter$count = 85807;
	#10 counter$count = 85808;
	#10 counter$count = 85809;
	#10 counter$count = 85810;
	#10 counter$count = 85811;
	#10 counter$count = 85812;
	#10 counter$count = 85813;
	#10 counter$count = 85814;
	#10 counter$count = 85815;
	#10 counter$count = 85816;
	#10 counter$count = 85817;
	#10 counter$count = 85818;
	#10 counter$count = 85819;
	#10 counter$count = 85820;
	#10 counter$count = 85821;
	#10 counter$count = 85822;
	#10 counter$count = 85823;
	#10 counter$count = 85824;
	#10 counter$count = 85825;
	#10 counter$count = 85826;
	#10 counter$count = 85827;
	#10 counter$count = 85828;
	#10 counter$count = 85829;
	#10 counter$count = 85830;
	#10 counter$count = 85831;
	#10 counter$count = 85832;
	#10 counter$count = 85833;
	#10 counter$count = 85834;
	#10 counter$count = 85835;
	#10 counter$count = 85836;
	#10 counter$count = 85837;
	#10 counter$count = 85838;
	#10 counter$count = 85839;
	#10 counter$count = 85840;
	#10 counter$count = 85841;
	#10 counter$count = 85842;
	#10 counter$count = 85843;
	#10 counter$count = 85844;
	#10 counter$count = 85845;
	#10 counter$count = 85846;
	#10 counter$count = 85847;
	#10 counter$count = 85848;
	#10 counter$count = 85849;
	#10 counter$count = 85850;
	#10 counter$count = 85851;
	#10 counter$count = 85852;
	#10 counter$count = 85853;
	#10 counter$count = 85854;
	#10 counter$count = 85855;
	#10 counter$count = 85856;
	#10 counter$count = 85857;
	#10 counter$count = 85858;
	#10 counter$count = 85859;
	#10 counter$count = 85860;
	#10 counter$count = 85861;
	#10 counter$count = 85862;
	#10 counter$count = 85863;
	#10 counter$count = 85864;
	#10 counter$count = 85865;
	#10 counter$count = 85866;
	#10 counter$count = 85867;
	#10 counter$count = 85868;
	#10 counter$count = 85869;
	#10 counter$count = 85870;
	#10 counter$count = 85871;
	#10 counter$count = 85872;
	#10 counter$count = 85873;
	#10 counter$count = 85874;
	#10 counter$count = 85875;
	#10 counter$count = 85876;
	#10 counter$count = 85877;
	#10 counter$count = 85878;
	#10 counter$count = 85879;
	#10 counter$count = 85880;
	#10 counter$count = 85881;
	#10 counter$count = 85882;
	#10 counter$count = 85883;
	#10 counter$count = 85884;
	#10 counter$count = 85885;
	#10 counter$count = 85886;
	#10 counter$count = 85887;
	#10 counter$count = 85888;
	#10 counter$count = 85889;
	#10 counter$count = 85890;
	#10 counter$count = 85891;
	#10 counter$count = 85892;
	#10 counter$count = 85893;
	#10 counter$count = 85894;
	#10 counter$count = 85895;
	#10 counter$count = 85896;
	#10 counter$count = 85897;
	#10 counter$count = 85898;
	#10 counter$count = 85899;
	#10 counter$count = 85900;
	#10 counter$count = 85901;
	#10 counter$count = 85902;
	#10 counter$count = 85903;
	#10 counter$count = 85904;
	#10 counter$count = 85905;
	#10 counter$count = 85906;
	#10 counter$count = 85907;
	#10 counter$count = 85908;
	#10 counter$count = 85909;
	#10 counter$count = 85910;
	#10 counter$count = 85911;
	#10 counter$count = 85912;
	#10 counter$count = 85913;
	#10 counter$count = 85914;
	#10 counter$count = 85915;
	#10 counter$count = 85916;
	#10 counter$count = 85917;
	#10 counter$count = 85918;
	#10 counter$count = 85919;
	#10 counter$count = 85920;
	#10 counter$count = 85921;
	#10 counter$count = 85922;
	#10 counter$count = 85923;
	#10 counter$count = 85924;
	#10 counter$count = 85925;
	#10 counter$count = 85926;
	#10 counter$count = 85927;
	#10 counter$count = 85928;
	#10 counter$count = 85929;
	#10 counter$count = 85930;
	#10 counter$count = 85931;
	#10 counter$count = 85932;
	#10 counter$count = 85933;
	#10 counter$count = 85934;
	#10 counter$count = 85935;
	#10 counter$count = 85936;
	#10 counter$count = 85937;
	#10 counter$count = 85938;
	#10 counter$count = 85939;
	#10 counter$count = 85940;
	#10 counter$count = 85941;
	#10 counter$count = 85942;
	#10 counter$count = 85943;
	#10 counter$count = 85944;
	#10 counter$count = 85945;
	#10 counter$count = 85946;
	#10 counter$count = 85947;
	#10 counter$count = 85948;
	#10 counter$count = 85949;
	#10 counter$count = 85950;
	#10 counter$count = 85951;
	#10 counter$count = 85952;
	#10 counter$count = 85953;
	#10 counter$count = 85954;
	#10 counter$count = 85955;
	#10 counter$count = 85956;
	#10 counter$count = 85957;
	#10 counter$count = 85958;
	#10 counter$count = 85959;
	#10 counter$count = 85960;
	#10 counter$count = 85961;
	#10 counter$count = 85962;
	#10 counter$count = 85963;
	#10 counter$count = 85964;
	#10 counter$count = 85965;
	#10 counter$count = 85966;
	#10 counter$count = 85967;
	#10 counter$count = 85968;
	#10 counter$count = 85969;
	#10 counter$count = 85970;
	#10 counter$count = 85971;
	#10 counter$count = 85972;
	#10 counter$count = 85973;
	#10 counter$count = 85974;
	#10 counter$count = 85975;
	#10 counter$count = 85976;
	#10 counter$count = 85977;
	#10 counter$count = 85978;
	#10 counter$count = 85979;
	#10 counter$count = 85980;
	#10 counter$count = 85981;
	#10 counter$count = 85982;
	#10 counter$count = 85983;
	#10 counter$count = 85984;
	#10 counter$count = 85985;
	#10 counter$count = 85986;
	#10 counter$count = 85987;
	#10 counter$count = 85988;
	#10 counter$count = 85989;
	#10 counter$count = 85990;
	#10 counter$count = 85991;
	#10 counter$count = 85992;
	#10 counter$count = 85993;
	#10 counter$count = 85994;
	#10 counter$count = 85995;
	#10 counter$count = 85996;
	#10 counter$count = 85997;
	#10 counter$count = 85998;
	#10 counter$count = 85999;
	#10 counter$count = 86000;
	#10 counter$count = 86001;
	#10 counter$count = 86002;
	#10 counter$count = 86003;
	#10 counter$count = 86004;
	#10 counter$count = 86005;
	#10 counter$count = 86006;
	#10 counter$count = 86007;
	#10 counter$count = 86008;
	#10 counter$count = 86009;
	#10 counter$count = 86010;
	#10 counter$count = 86011;
	#10 counter$count = 86012;
	#10 counter$count = 86013;
	#10 counter$count = 86014;
	#10 counter$count = 86015;
	#10 counter$count = 86016;
	#10 counter$count = 86017;
	#10 counter$count = 86018;
	#10 counter$count = 86019;
	#10 counter$count = 86020;
	#10 counter$count = 86021;
	#10 counter$count = 86022;
	#10 counter$count = 86023;
	#10 counter$count = 86024;
	#10 counter$count = 86025;
	#10 counter$count = 86026;
	#10 counter$count = 86027;
	#10 counter$count = 86028;
	#10 counter$count = 86029;
	#10 counter$count = 86030;
	#10 counter$count = 86031;
	#10 counter$count = 86032;
	#10 counter$count = 86033;
	#10 counter$count = 86034;
	#10 counter$count = 86035;
	#10 counter$count = 86036;
	#10 counter$count = 86037;
	#10 counter$count = 86038;
	#10 counter$count = 86039;
	#10 counter$count = 86040;
	#10 counter$count = 86041;
	#10 counter$count = 86042;
	#10 counter$count = 86043;
	#10 counter$count = 86044;
	#10 counter$count = 86045;
	#10 counter$count = 86046;
	#10 counter$count = 86047;
	#10 counter$count = 86048;
	#10 counter$count = 86049;
	#10 counter$count = 86050;
	#10 counter$count = 86051;
	#10 counter$count = 86052;
	#10 counter$count = 86053;
	#10 counter$count = 86054;
	#10 counter$count = 86055;
	#10 counter$count = 86056;
	#10 counter$count = 86057;
	#10 counter$count = 86058;
	#10 counter$count = 86059;
	#10 counter$count = 86060;
	#10 counter$count = 86061;
	#10 counter$count = 86062;
	#10 counter$count = 86063;
	#10 counter$count = 86064;
	#10 counter$count = 86065;
	#10 counter$count = 86066;
	#10 counter$count = 86067;
	#10 counter$count = 86068;
	#10 counter$count = 86069;
	#10 counter$count = 86070;
	#10 counter$count = 86071;
	#10 counter$count = 86072;
	#10 counter$count = 86073;
	#10 counter$count = 86074;
	#10 counter$count = 86075;
	#10 counter$count = 86076;
	#10 counter$count = 86077;
	#10 counter$count = 86078;
	#10 counter$count = 86079;
	#10 counter$count = 86080;
	#10 counter$count = 86081;
	#10 counter$count = 86082;
	#10 counter$count = 86083;
	#10 counter$count = 86084;
	#10 counter$count = 86085;
	#10 counter$count = 86086;
	#10 counter$count = 86087;
	#10 counter$count = 86088;
	#10 counter$count = 86089;
	#10 counter$count = 86090;
	#10 counter$count = 86091;
	#10 counter$count = 86092;
	#10 counter$count = 86093;
	#10 counter$count = 86094;
	#10 counter$count = 86095;
	#10 counter$count = 86096;
	#10 counter$count = 86097;
	#10 counter$count = 86098;
	#10 counter$count = 86099;
	#10 counter$count = 86100;
	#10 counter$count = 86101;
	#10 counter$count = 86102;
	#10 counter$count = 86103;
	#10 counter$count = 86104;
	#10 counter$count = 86105;
	#10 counter$count = 86106;
	#10 counter$count = 86107;
	#10 counter$count = 86108;
	#10 counter$count = 86109;
	#10 counter$count = 86110;
	#10 counter$count = 86111;
	#10 counter$count = 86112;
	#10 counter$count = 86113;
	#10 counter$count = 86114;
	#10 counter$count = 86115;
	#10 counter$count = 86116;
	#10 counter$count = 86117;
	#10 counter$count = 86118;
	#10 counter$count = 86119;
	#10 counter$count = 86120;
	#10 counter$count = 86121;
	#10 counter$count = 86122;
	#10 counter$count = 86123;
	#10 counter$count = 86124;
	#10 counter$count = 86125;
	#10 counter$count = 86126;
	#10 counter$count = 86127;
	#10 counter$count = 86128;
	#10 counter$count = 86129;
	#10 counter$count = 86130;
	#10 counter$count = 86131;
	#10 counter$count = 86132;
	#10 counter$count = 86133;
	#10 counter$count = 86134;
	#10 counter$count = 86135;
	#10 counter$count = 86136;
	#10 counter$count = 86137;
	#10 counter$count = 86138;
	#10 counter$count = 86139;
	#10 counter$count = 86140;
	#10 counter$count = 86141;
	#10 counter$count = 86142;
	#10 counter$count = 86143;
	#10 counter$count = 86144;
	#10 counter$count = 86145;
	#10 counter$count = 86146;
	#10 counter$count = 86147;
	#10 counter$count = 86148;
	#10 counter$count = 86149;
	#10 counter$count = 86150;
	#10 counter$count = 86151;
	#10 counter$count = 86152;
	#10 counter$count = 86153;
	#10 counter$count = 86154;
	#10 counter$count = 86155;
	#10 counter$count = 86156;
	#10 counter$count = 86157;
	#10 counter$count = 86158;
	#10 counter$count = 86159;
	#10 counter$count = 86160;
	#10 counter$count = 86161;
	#10 counter$count = 86162;
	#10 counter$count = 86163;
	#10 counter$count = 86164;
	#10 counter$count = 86165;
	#10 counter$count = 86166;
	#10 counter$count = 86167;
	#10 counter$count = 86168;
	#10 counter$count = 86169;
	#10 counter$count = 86170;
	#10 counter$count = 86171;
	#10 counter$count = 86172;
	#10 counter$count = 86173;
	#10 counter$count = 86174;
	#10 counter$count = 86175;
	#10 counter$count = 86176;
	#10 counter$count = 86177;
	#10 counter$count = 86178;
	#10 counter$count = 86179;
	#10 counter$count = 86180;
	#10 counter$count = 86181;
	#10 counter$count = 86182;
	#10 counter$count = 86183;
	#10 counter$count = 86184;
	#10 counter$count = 86185;
	#10 counter$count = 86186;
	#10 counter$count = 86187;
	#10 counter$count = 86188;
	#10 counter$count = 86189;
	#10 counter$count = 86190;
	#10 counter$count = 86191;
	#10 counter$count = 86192;
	#10 counter$count = 86193;
	#10 counter$count = 86194;
	#10 counter$count = 86195;
	#10 counter$count = 86196;
	#10 counter$count = 86197;
	#10 counter$count = 86198;
	#10 counter$count = 86199;
	#10 counter$count = 86200;
	#10 counter$count = 86201;
	#10 counter$count = 86202;
	#10 counter$count = 86203;
	#10 counter$count = 86204;
	#10 counter$count = 86205;
	#10 counter$count = 86206;
	#10 counter$count = 86207;
	#10 counter$count = 86208;
	#10 counter$count = 86209;
	#10 counter$count = 86210;
	#10 counter$count = 86211;
	#10 counter$count = 86212;
	#10 counter$count = 86213;
	#10 counter$count = 86214;
	#10 counter$count = 86215;
	#10 counter$count = 86216;
	#10 counter$count = 86217;
	#10 counter$count = 86218;
	#10 counter$count = 86219;
	#10 counter$count = 86220;
	#10 counter$count = 86221;
	#10 counter$count = 86222;
	#10 counter$count = 86223;
	#10 counter$count = 86224;
	#10 counter$count = 86225;
	#10 counter$count = 86226;
	#10 counter$count = 86227;
	#10 counter$count = 86228;
	#10 counter$count = 86229;
	#10 counter$count = 86230;
	#10 counter$count = 86231;
	#10 counter$count = 86232;
	#10 counter$count = 86233;
	#10 counter$count = 86234;
	#10 counter$count = 86235;
	#10 counter$count = 86236;
	#10 counter$count = 86237;
	#10 counter$count = 86238;
	#10 counter$count = 86239;
	#10 counter$count = 86240;
	#10 counter$count = 86241;
	#10 counter$count = 86242;
	#10 counter$count = 86243;
	#10 counter$count = 86244;
	#10 counter$count = 86245;
	#10 counter$count = 86246;
	#10 counter$count = 86247;
	#10 counter$count = 86248;
	#10 counter$count = 86249;
	#10 counter$count = 86250;
	#10 counter$count = 86251;
	#10 counter$count = 86252;
	#10 counter$count = 86253;
	#10 counter$count = 86254;
	#10 counter$count = 86255;
	#10 counter$count = 86256;
	#10 counter$count = 86257;
	#10 counter$count = 86258;
	#10 counter$count = 86259;
	#10 counter$count = 86260;
	#10 counter$count = 86261;
	#10 counter$count = 86262;
	#10 counter$count = 86263;
	#10 counter$count = 86264;
	#10 counter$count = 86265;
	#10 counter$count = 86266;
	#10 counter$count = 86267;
	#10 counter$count = 86268;
	#10 counter$count = 86269;
	#10 counter$count = 86270;
	#10 counter$count = 86271;
	#10 counter$count = 86272;
	#10 counter$count = 86273;
	#10 counter$count = 86274;
	#10 counter$count = 86275;
	#10 counter$count = 86276;
	#10 counter$count = 86277;
	#10 counter$count = 86278;
	#10 counter$count = 86279;
	#10 counter$count = 86280;
	#10 counter$count = 86281;
	#10 counter$count = 86282;
	#10 counter$count = 86283;
	#10 counter$count = 86284;
	#10 counter$count = 86285;
	#10 counter$count = 86286;
	#10 counter$count = 86287;
	#10 counter$count = 86288;
	#10 counter$count = 86289;
	#10 counter$count = 86290;
	#10 counter$count = 86291;
	#10 counter$count = 86292;
	#10 counter$count = 86293;
	#10 counter$count = 86294;
	#10 counter$count = 86295;
	#10 counter$count = 86296;
	#10 counter$count = 86297;
	#10 counter$count = 86298;
	#10 counter$count = 86299;
	#10 counter$count = 86300;
	#10 counter$count = 86301;
	#10 counter$count = 86302;
	#10 counter$count = 86303;
	#10 counter$count = 86304;
	#10 counter$count = 86305;
	#10 counter$count = 86306;
	#10 counter$count = 86307;
	#10 counter$count = 86308;
	#10 counter$count = 86309;
	#10 counter$count = 86310;
	#10 counter$count = 86311;
	#10 counter$count = 86312;
	#10 counter$count = 86313;
	#10 counter$count = 86314;
	#10 counter$count = 86315;
	#10 counter$count = 86316;
	#10 counter$count = 86317;
	#10 counter$count = 86318;
	#10 counter$count = 86319;
	#10 counter$count = 86320;
	#10 counter$count = 86321;
	#10 counter$count = 86322;
	#10 counter$count = 86323;
	#10 counter$count = 86324;
	#10 counter$count = 86325;
	#10 counter$count = 86326;
	#10 counter$count = 86327;
	#10 counter$count = 86328;
	#10 counter$count = 86329;
	#10 counter$count = 86330;
	#10 counter$count = 86331;
	#10 counter$count = 86332;
	#10 counter$count = 86333;
	#10 counter$count = 86334;
	#10 counter$count = 86335;
	#10 counter$count = 86336;
	#10 counter$count = 86337;
	#10 counter$count = 86338;
	#10 counter$count = 86339;
	#10 counter$count = 86340;
	#10 counter$count = 86341;
	#10 counter$count = 86342;
	#10 counter$count = 86343;
	#10 counter$count = 86344;
	#10 counter$count = 86345;
	#10 counter$count = 86346;
	#10 counter$count = 86347;
	#10 counter$count = 86348;
	#10 counter$count = 86349;
	#10 counter$count = 86350;
	#10 counter$count = 86351;
	#10 counter$count = 86352;
	#10 counter$count = 86353;
	#10 counter$count = 86354;
	#10 counter$count = 86355;
	#10 counter$count = 86356;
	#10 counter$count = 86357;
	#10 counter$count = 86358;
	#10 counter$count = 86359;
	#10 counter$count = 86360;
	#10 counter$count = 86361;
	#10 counter$count = 86362;
	#10 counter$count = 86363;
	#10 counter$count = 86364;
	#10 counter$count = 86365;
	#10 counter$count = 86366;
	#10 counter$count = 86367;
	#10 counter$count = 86368;
	#10 counter$count = 86369;
	#10 counter$count = 86370;
	#10 counter$count = 86371;
	#10 counter$count = 86372;
	#10 counter$count = 86373;
	#10 counter$count = 86374;
	#10 counter$count = 86375;
	#10 counter$count = 86376;
	#10 counter$count = 86377;
	#10 counter$count = 86378;
	#10 counter$count = 86379;
	#10 counter$count = 86380;
	#10 counter$count = 86381;
	#10 counter$count = 86382;
	#10 counter$count = 86383;
	#10 counter$count = 86384;
	#10 counter$count = 86385;
	#10 counter$count = 86386;
	#10 counter$count = 86387;
	#10 counter$count = 86388;
	#10 counter$count = 86389;
	#10 counter$count = 86390;
	#10 counter$count = 86391;
	#10 counter$count = 86392;
	#10 counter$count = 86393;
	#10 counter$count = 86394;
	#10 counter$count = 86395;
	#10 counter$count = 86396;
	#10 counter$count = 86397;
	#10 counter$count = 86398;
	#10 counter$count = 86399;
	#10 counter$count = 86400;
	#10 counter$count = 86401;
	#10 counter$count = 86402;
	#10 counter$count = 86403;
	#10 counter$count = 86404;
	#10 counter$count = 86405;
	#10 counter$count = 86406;
	#10 counter$count = 86407;
	#10 counter$count = 86408;
	#10 counter$count = 86409;
	#10 counter$count = 86410;
	#10 counter$count = 86411;
	#10 counter$count = 86412;
	#10 counter$count = 86413;
	#10 counter$count = 86414;
	#10 counter$count = 86415;
	#10 counter$count = 86416;
	#10 counter$count = 86417;
	#10 counter$count = 86418;
	#10 counter$count = 86419;
	#10 counter$count = 86420;
	#10 counter$count = 86421;
	#10 counter$count = 86422;
	#10 counter$count = 86423;
	#10 counter$count = 86424;
	#10 counter$count = 86425;
	#10 counter$count = 86426;
	#10 counter$count = 86427;
	#10 counter$count = 86428;
	#10 counter$count = 86429;
	#10 counter$count = 86430;
	#10 counter$count = 86431;
	#10 counter$count = 86432;
	#10 counter$count = 86433;
	#10 counter$count = 86434;
	#10 counter$count = 86435;
	#10 counter$count = 86436;
	#10 counter$count = 86437;
	#10 counter$count = 86438;
	#10 counter$count = 86439;
	#10 counter$count = 86440;
	#10 counter$count = 86441;
	#10 counter$count = 86442;
	#10 counter$count = 86443;
	#10 counter$count = 86444;
	#10 counter$count = 86445;
	#10 counter$count = 86446;
	#10 counter$count = 86447;
	#10 counter$count = 86448;
	#10 counter$count = 86449;
	#10 counter$count = 86450;
	#10 counter$count = 86451;
	#10 counter$count = 86452;
	#10 counter$count = 86453;
	#10 counter$count = 86454;
	#10 counter$count = 86455;
	#10 counter$count = 86456;
	#10 counter$count = 86457;
	#10 counter$count = 86458;
	#10 counter$count = 86459;
	#10 counter$count = 86460;
	#10 counter$count = 86461;
	#10 counter$count = 86462;
	#10 counter$count = 86463;
	#10 counter$count = 86464;
	#10 counter$count = 86465;
	#10 counter$count = 86466;
	#10 counter$count = 86467;
	#10 counter$count = 86468;
	#10 counter$count = 86469;
	#10 counter$count = 86470;
	#10 counter$count = 86471;
	#10 counter$count = 86472;
	#10 counter$count = 86473;
	#10 counter$count = 86474;
	#10 counter$count = 86475;
	#10 counter$count = 86476;
	#10 counter$count = 86477;
	#10 counter$count = 86478;
	#10 counter$count = 86479;
	#10 counter$count = 86480;
	#10 counter$count = 86481;
	#10 counter$count = 86482;
	#10 counter$count = 86483;
	#10 counter$count = 86484;
	#10 counter$count = 86485;
	#10 counter$count = 86486;
	#10 counter$count = 86487;
	#10 counter$count = 86488;
	#10 counter$count = 86489;
	#10 counter$count = 86490;
	#10 counter$count = 86491;
	#10 counter$count = 86492;
	#10 counter$count = 86493;
	#10 counter$count = 86494;
	#10 counter$count = 86495;
	#10 counter$count = 86496;
	#10 counter$count = 86497;
	#10 counter$count = 86498;
	#10 counter$count = 86499;
	#10 counter$count = 86500;
	#10 counter$count = 86501;
	#10 counter$count = 86502;
	#10 counter$count = 86503;
	#10 counter$count = 86504;
	#10 counter$count = 86505;
	#10 counter$count = 86506;
	#10 counter$count = 86507;
	#10 counter$count = 86508;
	#10 counter$count = 86509;
	#10 counter$count = 86510;
	#10 counter$count = 86511;
	#10 counter$count = 86512;
	#10 counter$count = 86513;
	#10 counter$count = 86514;
	#10 counter$count = 86515;
	#10 counter$count = 86516;
	#10 counter$count = 86517;
	#10 counter$count = 86518;
	#10 counter$count = 86519;
	#10 counter$count = 86520;
	#10 counter$count = 86521;
	#10 counter$count = 86522;
	#10 counter$count = 86523;
	#10 counter$count = 86524;
	#10 counter$count = 86525;
	#10 counter$count = 86526;
	#10 counter$count = 86527;
	#10 counter$count = 86528;
	#10 counter$count = 86529;
	#10 counter$count = 86530;
	#10 counter$count = 86531;
	#10 counter$count = 86532;
	#10 counter$count = 86533;
	#10 counter$count = 86534;
	#10 counter$count = 86535;
	#10 counter$count = 86536;
	#10 counter$count = 86537;
	#10 counter$count = 86538;
	#10 counter$count = 86539;
	#10 counter$count = 86540;
	#10 counter$count = 86541;
	#10 counter$count = 86542;
	#10 counter$count = 86543;
	#10 counter$count = 86544;
	#10 counter$count = 86545;
	#10 counter$count = 86546;
	#10 counter$count = 86547;
	#10 counter$count = 86548;
	#10 counter$count = 86549;
	#10 counter$count = 86550;
	#10 counter$count = 86551;
	#10 counter$count = 86552;
	#10 counter$count = 86553;
	#10 counter$count = 86554;
	#10 counter$count = 86555;
	#10 counter$count = 86556;
	#10 counter$count = 86557;
	#10 counter$count = 86558;
	#10 counter$count = 86559;
	#10 counter$count = 86560;
	#10 counter$count = 86561;
	#10 counter$count = 86562;
	#10 counter$count = 86563;
	#10 counter$count = 86564;
	#10 counter$count = 86565;
	#10 counter$count = 86566;
	#10 counter$count = 86567;
	#10 counter$count = 86568;
	#10 counter$count = 86569;
	#10 counter$count = 86570;
	#10 counter$count = 86571;
	#10 counter$count = 86572;
	#10 counter$count = 86573;
	#10 counter$count = 86574;
	#10 counter$count = 86575;
	#10 counter$count = 86576;
	#10 counter$count = 86577;
	#10 counter$count = 86578;
	#10 counter$count = 86579;
	#10 counter$count = 86580;
	#10 counter$count = 86581;
	#10 counter$count = 86582;
	#10 counter$count = 86583;
	#10 counter$count = 86584;
	#10 counter$count = 86585;
	#10 counter$count = 86586;
	#10 counter$count = 86587;
	#10 counter$count = 86588;
	#10 counter$count = 86589;
	#10 counter$count = 86590;
	#10 counter$count = 86591;
	#10 counter$count = 86592;
	#10 counter$count = 86593;
	#10 counter$count = 86594;
	#10 counter$count = 86595;
	#10 counter$count = 86596;
	#10 counter$count = 86597;
	#10 counter$count = 86598;
	#10 counter$count = 86599;
	#10 counter$count = 86600;
	#10 counter$count = 86601;
	#10 counter$count = 86602;
	#10 counter$count = 86603;
	#10 counter$count = 86604;
	#10 counter$count = 86605;
	#10 counter$count = 86606;
	#10 counter$count = 86607;
	#10 counter$count = 86608;
	#10 counter$count = 86609;
	#10 counter$count = 86610;
	#10 counter$count = 86611;
	#10 counter$count = 86612;
	#10 counter$count = 86613;
	#10 counter$count = 86614;
	#10 counter$count = 86615;
	#10 counter$count = 86616;
	#10 counter$count = 86617;
	#10 counter$count = 86618;
	#10 counter$count = 86619;
	#10 counter$count = 86620;
	#10 counter$count = 86621;
	#10 counter$count = 86622;
	#10 counter$count = 86623;
	#10 counter$count = 86624;
	#10 counter$count = 86625;
	#10 counter$count = 86626;
	#10 counter$count = 86627;
	#10 counter$count = 86628;
	#10 counter$count = 86629;
	#10 counter$count = 86630;
	#10 counter$count = 86631;
	#10 counter$count = 86632;
	#10 counter$count = 86633;
	#10 counter$count = 86634;
	#10 counter$count = 86635;
	#10 counter$count = 86636;
	#10 counter$count = 86637;
	#10 counter$count = 86638;
	#10 counter$count = 86639;
	#10 counter$count = 86640;
	#10 counter$count = 86641;
	#10 counter$count = 86642;
	#10 counter$count = 86643;
	#10 counter$count = 86644;
	#10 counter$count = 86645;
	#10 counter$count = 86646;
	#10 counter$count = 86647;
	#10 counter$count = 86648;
	#10 counter$count = 86649;
	#10 counter$count = 86650;
	#10 counter$count = 86651;
	#10 counter$count = 86652;
	#10 counter$count = 86653;
	#10 counter$count = 86654;
	#10 counter$count = 86655;
	#10 counter$count = 86656;
	#10 counter$count = 86657;
	#10 counter$count = 86658;
	#10 counter$count = 86659;
	#10 counter$count = 86660;
	#10 counter$count = 86661;
	#10 counter$count = 86662;
	#10 counter$count = 86663;
	#10 counter$count = 86664;
	#10 counter$count = 86665;
	#10 counter$count = 86666;
	#10 counter$count = 86667;
	#10 counter$count = 86668;
	#10 counter$count = 86669;
	#10 counter$count = 86670;
	#10 counter$count = 86671;
	#10 counter$count = 86672;
	#10 counter$count = 86673;
	#10 counter$count = 86674;
	#10 counter$count = 86675;
	#10 counter$count = 86676;
	#10 counter$count = 86677;
	#10 counter$count = 86678;
	#10 counter$count = 86679;
	#10 counter$count = 86680;
	#10 counter$count = 86681;
	#10 counter$count = 86682;
	#10 counter$count = 86683;
	#10 counter$count = 86684;
	#10 counter$count = 86685;
	#10 counter$count = 86686;
	#10 counter$count = 86687;
	#10 counter$count = 86688;
	#10 counter$count = 86689;
	#10 counter$count = 86690;
	#10 counter$count = 86691;
	#10 counter$count = 86692;
	#10 counter$count = 86693;
	#10 counter$count = 86694;
	#10 counter$count = 86695;
	#10 counter$count = 86696;
	#10 counter$count = 86697;
	#10 counter$count = 86698;
	#10 counter$count = 86699;
	#10 counter$count = 86700;
	#10 counter$count = 86701;
	#10 counter$count = 86702;
	#10 counter$count = 86703;
	#10 counter$count = 86704;
	#10 counter$count = 86705;
	#10 counter$count = 86706;
	#10 counter$count = 86707;
	#10 counter$count = 86708;
	#10 counter$count = 86709;
	#10 counter$count = 86710;
	#10 counter$count = 86711;
	#10 counter$count = 86712;
	#10 counter$count = 86713;
	#10 counter$count = 86714;
	#10 counter$count = 86715;
	#10 counter$count = 86716;
	#10 counter$count = 86717;
	#10 counter$count = 86718;
	#10 counter$count = 86719;
	#10 counter$count = 86720;
	#10 counter$count = 86721;
	#10 counter$count = 86722;
	#10 counter$count = 86723;
	#10 counter$count = 86724;
	#10 counter$count = 86725;
	#10 counter$count = 86726;
	#10 counter$count = 86727;
	#10 counter$count = 86728;
	#10 counter$count = 86729;
	#10 counter$count = 86730;
	#10 counter$count = 86731;
	#10 counter$count = 86732;
	#10 counter$count = 86733;
	#10 counter$count = 86734;
	#10 counter$count = 86735;
	#10 counter$count = 86736;
	#10 counter$count = 86737;
	#10 counter$count = 86738;
	#10 counter$count = 86739;
	#10 counter$count = 86740;
	#10 counter$count = 86741;
	#10 counter$count = 86742;
	#10 counter$count = 86743;
	#10 counter$count = 86744;
	#10 counter$count = 86745;
	#10 counter$count = 86746;
	#10 counter$count = 86747;
	#10 counter$count = 86748;
	#10 counter$count = 86749;
	#10 counter$count = 86750;
	#10 counter$count = 86751;
	#10 counter$count = 86752;
	#10 counter$count = 86753;
	#10 counter$count = 86754;
	#10 counter$count = 86755;
	#10 counter$count = 86756;
	#10 counter$count = 86757;
	#10 counter$count = 86758;
	#10 counter$count = 86759;
	#10 counter$count = 86760;
	#10 counter$count = 86761;
	#10 counter$count = 86762;
	#10 counter$count = 86763;
	#10 counter$count = 86764;
	#10 counter$count = 86765;
	#10 counter$count = 86766;
	#10 counter$count = 86767;
	#10 counter$count = 86768;
	#10 counter$count = 86769;
	#10 counter$count = 86770;
	#10 counter$count = 86771;
	#10 counter$count = 86772;
	#10 counter$count = 86773;
	#10 counter$count = 86774;
	#10 counter$count = 86775;
	#10 counter$count = 86776;
	#10 counter$count = 86777;
	#10 counter$count = 86778;
	#10 counter$count = 86779;
	#10 counter$count = 86780;
	#10 counter$count = 86781;
	#10 counter$count = 86782;
	#10 counter$count = 86783;
	#10 counter$count = 86784;
	#10 counter$count = 86785;
	#10 counter$count = 86786;
	#10 counter$count = 86787;
	#10 counter$count = 86788;
	#10 counter$count = 86789;
	#10 counter$count = 86790;
	#10 counter$count = 86791;
	#10 counter$count = 86792;
	#10 counter$count = 86793;
	#10 counter$count = 86794;
	#10 counter$count = 86795;
	#10 counter$count = 86796;
	#10 counter$count = 86797;
	#10 counter$count = 86798;
	#10 counter$count = 86799;
	#10 counter$count = 86800;
	#10 counter$count = 86801;
	#10 counter$count = 86802;
	#10 counter$count = 86803;
	#10 counter$count = 86804;
	#10 counter$count = 86805;
	#10 counter$count = 86806;
	#10 counter$count = 86807;
	#10 counter$count = 86808;
	#10 counter$count = 86809;
	#10 counter$count = 86810;
	#10 counter$count = 86811;
	#10 counter$count = 86812;
	#10 counter$count = 86813;
	#10 counter$count = 86814;
	#10 counter$count = 86815;
	#10 counter$count = 86816;
	#10 counter$count = 86817;
	#10 counter$count = 86818;
	#10 counter$count = 86819;
	#10 counter$count = 86820;
	#10 counter$count = 86821;
	#10 counter$count = 86822;
	#10 counter$count = 86823;
	#10 counter$count = 86824;
	#10 counter$count = 86825;
	#10 counter$count = 86826;
	#10 counter$count = 86827;
	#10 counter$count = 86828;
	#10 counter$count = 86829;
	#10 counter$count = 86830;
	#10 counter$count = 86831;
	#10 counter$count = 86832;
	#10 counter$count = 86833;
	#10 counter$count = 86834;
	#10 counter$count = 86835;
	#10 counter$count = 86836;
	#10 counter$count = 86837;
	#10 counter$count = 86838;
	#10 counter$count = 86839;
	#10 counter$count = 86840;
	#10 counter$count = 86841;
	#10 counter$count = 86842;
	#10 counter$count = 86843;
	#10 counter$count = 86844;
	#10 counter$count = 86845;
	#10 counter$count = 86846;
	#10 counter$count = 86847;
	#10 counter$count = 86848;
	#10 counter$count = 86849;
	#10 counter$count = 86850;
	#10 counter$count = 86851;
	#10 counter$count = 86852;
	#10 counter$count = 86853;
	#10 counter$count = 86854;
	#10 counter$count = 86855;
	#10 counter$count = 86856;
	#10 counter$count = 86857;
	#10 counter$count = 86858;
	#10 counter$count = 86859;
	#10 counter$count = 86860;
	#10 counter$count = 86861;
	#10 counter$count = 86862;
	#10 counter$count = 86863;
	#10 counter$count = 86864;
	#10 counter$count = 86865;
	#10 counter$count = 86866;
	#10 counter$count = 86867;
	#10 counter$count = 86868;
	#10 counter$count = 86869;
	#10 counter$count = 86870;
	#10 counter$count = 86871;
	#10 counter$count = 86872;
	#10 counter$count = 86873;
	#10 counter$count = 86874;
	#10 counter$count = 86875;
	#10 counter$count = 86876;
	#10 counter$count = 86877;
	#10 counter$count = 86878;
	#10 counter$count = 86879;
	#10 counter$count = 86880;
	#10 counter$count = 86881;
	#10 counter$count = 86882;
	#10 counter$count = 86883;
	#10 counter$count = 86884;
	#10 counter$count = 86885;
	#10 counter$count = 86886;
	#10 counter$count = 86887;
	#10 counter$count = 86888;
	#10 counter$count = 86889;
	#10 counter$count = 86890;
	#10 counter$count = 86891;
	#10 counter$count = 86892;
	#10 counter$count = 86893;
	#10 counter$count = 86894;
	#10 counter$count = 86895;
	#10 counter$count = 86896;
	#10 counter$count = 86897;
	#10 counter$count = 86898;
	#10 counter$count = 86899;
	#10 counter$count = 86900;
	#10 counter$count = 86901;
	#10 counter$count = 86902;
	#10 counter$count = 86903;
	#10 counter$count = 86904;
	#10 counter$count = 86905;
	#10 counter$count = 86906;
	#10 counter$count = 86907;
	#10 counter$count = 86908;
	#10 counter$count = 86909;
	#10 counter$count = 86910;
	#10 counter$count = 86911;
	#10 counter$count = 86912;
	#10 counter$count = 86913;
	#10 counter$count = 86914;
	#10 counter$count = 86915;
	#10 counter$count = 86916;
	#10 counter$count = 86917;
	#10 counter$count = 86918;
	#10 counter$count = 86919;
	#10 counter$count = 86920;
	#10 counter$count = 86921;
	#10 counter$count = 86922;
	#10 counter$count = 86923;
	#10 counter$count = 86924;
	#10 counter$count = 86925;
	#10 counter$count = 86926;
	#10 counter$count = 86927;
	#10 counter$count = 86928;
	#10 counter$count = 86929;
	#10 counter$count = 86930;
	#10 counter$count = 86931;
	#10 counter$count = 86932;
	#10 counter$count = 86933;
	#10 counter$count = 86934;
	#10 counter$count = 86935;
	#10 counter$count = 86936;
	#10 counter$count = 86937;
	#10 counter$count = 86938;
	#10 counter$count = 86939;
	#10 counter$count = 86940;
	#10 counter$count = 86941;
	#10 counter$count = 86942;
	#10 counter$count = 86943;
	#10 counter$count = 86944;
	#10 counter$count = 86945;
	#10 counter$count = 86946;
	#10 counter$count = 86947;
	#10 counter$count = 86948;
	#10 counter$count = 86949;
	#10 counter$count = 86950;
	#10 counter$count = 86951;
	#10 counter$count = 86952;
	#10 counter$count = 86953;
	#10 counter$count = 86954;
	#10 counter$count = 86955;
	#10 counter$count = 86956;
	#10 counter$count = 86957;
	#10 counter$count = 86958;
	#10 counter$count = 86959;
	#10 counter$count = 86960;
	#10 counter$count = 86961;
	#10 counter$count = 86962;
	#10 counter$count = 86963;
	#10 counter$count = 86964;
	#10 counter$count = 86965;
	#10 counter$count = 86966;
	#10 counter$count = 86967;
	#10 counter$count = 86968;
	#10 counter$count = 86969;
	#10 counter$count = 86970;
	#10 counter$count = 86971;
	#10 counter$count = 86972;
	#10 counter$count = 86973;
	#10 counter$count = 86974;
	#10 counter$count = 86975;
	#10 counter$count = 86976;
	#10 counter$count = 86977;
	#10 counter$count = 86978;
	#10 counter$count = 86979;
	#10 counter$count = 86980;
	#10 counter$count = 86981;
	#10 counter$count = 86982;
	#10 counter$count = 86983;
	#10 counter$count = 86984;
	#10 counter$count = 86985;
	#10 counter$count = 86986;
	#10 counter$count = 86987;
	#10 counter$count = 86988;
	#10 counter$count = 86989;
	#10 counter$count = 86990;
	#10 counter$count = 86991;
	#10 counter$count = 86992;
	#10 counter$count = 86993;
	#10 counter$count = 86994;
	#10 counter$count = 86995;
	#10 counter$count = 86996;
	#10 counter$count = 86997;
	#10 counter$count = 86998;
	#10 counter$count = 86999;
	#10 counter$count = 87000;
	#10 counter$count = 87001;
	#10 counter$count = 87002;
	#10 counter$count = 87003;
	#10 counter$count = 87004;
	#10 counter$count = 87005;
	#10 counter$count = 87006;
	#10 counter$count = 87007;
	#10 counter$count = 87008;
	#10 counter$count = 87009;
	#10 counter$count = 87010;
	#10 counter$count = 87011;
	#10 counter$count = 87012;
	#10 counter$count = 87013;
	#10 counter$count = 87014;
	#10 counter$count = 87015;
	#10 counter$count = 87016;
	#10 counter$count = 87017;
	#10 counter$count = 87018;
	#10 counter$count = 87019;
	#10 counter$count = 87020;
	#10 counter$count = 87021;
	#10 counter$count = 87022;
	#10 counter$count = 87023;
	#10 counter$count = 87024;
	#10 counter$count = 87025;
	#10 counter$count = 87026;
	#10 counter$count = 87027;
	#10 counter$count = 87028;
	#10 counter$count = 87029;
	#10 counter$count = 87030;
	#10 counter$count = 87031;
	#10 counter$count = 87032;
	#10 counter$count = 87033;
	#10 counter$count = 87034;
	#10 counter$count = 87035;
	#10 counter$count = 87036;
	#10 counter$count = 87037;
	#10 counter$count = 87038;
	#10 counter$count = 87039;
	#10 counter$count = 87040;
	#10 counter$count = 87041;
	#10 counter$count = 87042;
	#10 counter$count = 87043;
	#10 counter$count = 87044;
	#10 counter$count = 87045;
	#10 counter$count = 87046;
	#10 counter$count = 87047;
	#10 counter$count = 87048;
	#10 counter$count = 87049;
	#10 counter$count = 87050;
	#10 counter$count = 87051;
	#10 counter$count = 87052;
	#10 counter$count = 87053;
	#10 counter$count = 87054;
	#10 counter$count = 87055;
	#10 counter$count = 87056;
	#10 counter$count = 87057;
	#10 counter$count = 87058;
	#10 counter$count = 87059;
	#10 counter$count = 87060;
	#10 counter$count = 87061;
	#10 counter$count = 87062;
	#10 counter$count = 87063;
	#10 counter$count = 87064;
	#10 counter$count = 87065;
	#10 counter$count = 87066;
	#10 counter$count = 87067;
	#10 counter$count = 87068;
	#10 counter$count = 87069;
	#10 counter$count = 87070;
	#10 counter$count = 87071;
	#10 counter$count = 87072;
	#10 counter$count = 87073;
	#10 counter$count = 87074;
	#10 counter$count = 87075;
	#10 counter$count = 87076;
	#10 counter$count = 87077;
	#10 counter$count = 87078;
	#10 counter$count = 87079;
	#10 counter$count = 87080;
	#10 counter$count = 87081;
	#10 counter$count = 87082;
	#10 counter$count = 87083;
	#10 counter$count = 87084;
	#10 counter$count = 87085;
	#10 counter$count = 87086;
	#10 counter$count = 87087;
	#10 counter$count = 87088;
	#10 counter$count = 87089;
	#10 counter$count = 87090;
	#10 counter$count = 87091;
	#10 counter$count = 87092;
	#10 counter$count = 87093;
	#10 counter$count = 87094;
	#10 counter$count = 87095;
	#10 counter$count = 87096;
	#10 counter$count = 87097;
	#10 counter$count = 87098;
	#10 counter$count = 87099;
	#10 counter$count = 87100;
	#10 counter$count = 87101;
	#10 counter$count = 87102;
	#10 counter$count = 87103;
	#10 counter$count = 87104;
	#10 counter$count = 87105;
	#10 counter$count = 87106;
	#10 counter$count = 87107;
	#10 counter$count = 87108;
	#10 counter$count = 87109;
	#10 counter$count = 87110;
	#10 counter$count = 87111;
	#10 counter$count = 87112;
	#10 counter$count = 87113;
	#10 counter$count = 87114;
	#10 counter$count = 87115;
	#10 counter$count = 87116;
	#10 counter$count = 87117;
	#10 counter$count = 87118;
	#10 counter$count = 87119;
	#10 counter$count = 87120;
	#10 counter$count = 87121;
	#10 counter$count = 87122;
	#10 counter$count = 87123;
	#10 counter$count = 87124;
	#10 counter$count = 87125;
	#10 counter$count = 87126;
	#10 counter$count = 87127;
	#10 counter$count = 87128;
	#10 counter$count = 87129;
	#10 counter$count = 87130;
	#10 counter$count = 87131;
	#10 counter$count = 87132;
	#10 counter$count = 87133;
	#10 counter$count = 87134;
	#10 counter$count = 87135;
	#10 counter$count = 87136;
	#10 counter$count = 87137;
	#10 counter$count = 87138;
	#10 counter$count = 87139;
	#10 counter$count = 87140;
	#10 counter$count = 87141;
	#10 counter$count = 87142;
	#10 counter$count = 87143;
	#10 counter$count = 87144;
	#10 counter$count = 87145;
	#10 counter$count = 87146;
	#10 counter$count = 87147;
	#10 counter$count = 87148;
	#10 counter$count = 87149;
	#10 counter$count = 87150;
	#10 counter$count = 87151;
	#10 counter$count = 87152;
	#10 counter$count = 87153;
	#10 counter$count = 87154;
	#10 counter$count = 87155;
	#10 counter$count = 87156;
	#10 counter$count = 87157;
	#10 counter$count = 87158;
	#10 counter$count = 87159;
	#10 counter$count = 87160;
	#10 counter$count = 87161;
	#10 counter$count = 87162;
	#10 counter$count = 87163;
	#10 counter$count = 87164;
	#10 counter$count = 87165;
	#10 counter$count = 87166;
	#10 counter$count = 87167;
	#10 counter$count = 87168;
	#10 counter$count = 87169;
	#10 counter$count = 87170;
	#10 counter$count = 87171;
	#10 counter$count = 87172;
	#10 counter$count = 87173;
	#10 counter$count = 87174;
	#10 counter$count = 87175;
	#10 counter$count = 87176;
	#10 counter$count = 87177;
	#10 counter$count = 87178;
	#10 counter$count = 87179;
	#10 counter$count = 87180;
	#10 counter$count = 87181;
	#10 counter$count = 87182;
	#10 counter$count = 87183;
	#10 counter$count = 87184;
	#10 counter$count = 87185;
	#10 counter$count = 87186;
	#10 counter$count = 87187;
	#10 counter$count = 87188;
	#10 counter$count = 87189;
	#10 counter$count = 87190;
	#10 counter$count = 87191;
	#10 counter$count = 87192;
	#10 counter$count = 87193;
	#10 counter$count = 87194;
	#10 counter$count = 87195;
	#10 counter$count = 87196;
	#10 counter$count = 87197;
	#10 counter$count = 87198;
	#10 counter$count = 87199;
	#10 counter$count = 87200;
	#10 counter$count = 87201;
	#10 counter$count = 87202;
	#10 counter$count = 87203;
	#10 counter$count = 87204;
	#10 counter$count = 87205;
	#10 counter$count = 87206;
	#10 counter$count = 87207;
	#10 counter$count = 87208;
	#10 counter$count = 87209;
	#10 counter$count = 87210;
	#10 counter$count = 87211;
	#10 counter$count = 87212;
	#10 counter$count = 87213;
	#10 counter$count = 87214;
	#10 counter$count = 87215;
	#10 counter$count = 87216;
	#10 counter$count = 87217;
	#10 counter$count = 87218;
	#10 counter$count = 87219;
	#10 counter$count = 87220;
	#10 counter$count = 87221;
	#10 counter$count = 87222;
	#10 counter$count = 87223;
	#10 counter$count = 87224;
	#10 counter$count = 87225;
	#10 counter$count = 87226;
	#10 counter$count = 87227;
	#10 counter$count = 87228;
	#10 counter$count = 87229;
	#10 counter$count = 87230;
	#10 counter$count = 87231;
	#10 counter$count = 87232;
	#10 counter$count = 87233;
	#10 counter$count = 87234;
	#10 counter$count = 87235;
	#10 counter$count = 87236;
	#10 counter$count = 87237;
	#10 counter$count = 87238;
	#10 counter$count = 87239;
	#10 counter$count = 87240;
	#10 counter$count = 87241;
	#10 counter$count = 87242;
	#10 counter$count = 87243;
	#10 counter$count = 87244;
	#10 counter$count = 87245;
	#10 counter$count = 87246;
	#10 counter$count = 87247;
	#10 counter$count = 87248;
	#10 counter$count = 87249;
	#10 counter$count = 87250;
	#10 counter$count = 87251;
	#10 counter$count = 87252;
	#10 counter$count = 87253;
	#10 counter$count = 87254;
	#10 counter$count = 87255;
	#10 counter$count = 87256;
	#10 counter$count = 87257;
	#10 counter$count = 87258;
	#10 counter$count = 87259;
	#10 counter$count = 87260;
	#10 counter$count = 87261;
	#10 counter$count = 87262;
	#10 counter$count = 87263;
	#10 counter$count = 87264;
	#10 counter$count = 87265;
	#10 counter$count = 87266;
	#10 counter$count = 87267;
	#10 counter$count = 87268;
	#10 counter$count = 87269;
	#10 counter$count = 87270;
	#10 counter$count = 87271;
	#10 counter$count = 87272;
	#10 counter$count = 87273;
	#10 counter$count = 87274;
	#10 counter$count = 87275;
	#10 counter$count = 87276;
	#10 counter$count = 87277;
	#10 counter$count = 87278;
	#10 counter$count = 87279;
	#10 counter$count = 87280;
	#10 counter$count = 87281;
	#10 counter$count = 87282;
	#10 counter$count = 87283;
	#10 counter$count = 87284;
	#10 counter$count = 87285;
	#10 counter$count = 87286;
	#10 counter$count = 87287;
	#10 counter$count = 87288;
	#10 counter$count = 87289;
	#10 counter$count = 87290;
	#10 counter$count = 87291;
	#10 counter$count = 87292;
	#10 counter$count = 87293;
	#10 counter$count = 87294;
	#10 counter$count = 87295;
	#10 counter$count = 87296;
	#10 counter$count = 87297;
	#10 counter$count = 87298;
	#10 counter$count = 87299;
	#10 counter$count = 87300;
	#10 counter$count = 87301;
	#10 counter$count = 87302;
	#10 counter$count = 87303;
	#10 counter$count = 87304;
	#10 counter$count = 87305;
	#10 counter$count = 87306;
	#10 counter$count = 87307;
	#10 counter$count = 87308;
	#10 counter$count = 87309;
	#10 counter$count = 87310;
	#10 counter$count = 87311;
	#10 counter$count = 87312;
	#10 counter$count = 87313;
	#10 counter$count = 87314;
	#10 counter$count = 87315;
	#10 counter$count = 87316;
	#10 counter$count = 87317;
	#10 counter$count = 87318;
	#10 counter$count = 87319;
	#10 counter$count = 87320;
	#10 counter$count = 87321;
	#10 counter$count = 87322;
	#10 counter$count = 87323;
	#10 counter$count = 87324;
	#10 counter$count = 87325;
	#10 counter$count = 87326;
	#10 counter$count = 87327;
	#10 counter$count = 87328;
	#10 counter$count = 87329;
	#10 counter$count = 87330;
	#10 counter$count = 87331;
	#10 counter$count = 87332;
	#10 counter$count = 87333;
	#10 counter$count = 87334;
	#10 counter$count = 87335;
	#10 counter$count = 87336;
	#10 counter$count = 87337;
	#10 counter$count = 87338;
	#10 counter$count = 87339;
	#10 counter$count = 87340;
	#10 counter$count = 87341;
	#10 counter$count = 87342;
	#10 counter$count = 87343;
	#10 counter$count = 87344;
	#10 counter$count = 87345;
	#10 counter$count = 87346;
	#10 counter$count = 87347;
	#10 counter$count = 87348;
	#10 counter$count = 87349;
	#10 counter$count = 87350;
	#10 counter$count = 87351;
	#10 counter$count = 87352;
	#10 counter$count = 87353;
	#10 counter$count = 87354;
	#10 counter$count = 87355;
	#10 counter$count = 87356;
	#10 counter$count = 87357;
	#10 counter$count = 87358;
	#10 counter$count = 87359;
	#10 counter$count = 87360;
	#10 counter$count = 87361;
	#10 counter$count = 87362;
	#10 counter$count = 87363;
	#10 counter$count = 87364;
	#10 counter$count = 87365;
	#10 counter$count = 87366;
	#10 counter$count = 87367;
	#10 counter$count = 87368;
	#10 counter$count = 87369;
	#10 counter$count = 87370;
	#10 counter$count = 87371;
	#10 counter$count = 87372;
	#10 counter$count = 87373;
	#10 counter$count = 87374;
	#10 counter$count = 87375;
	#10 counter$count = 87376;
	#10 counter$count = 87377;
	#10 counter$count = 87378;
	#10 counter$count = 87379;
	#10 counter$count = 87380;
	#10 counter$count = 87381;
	#10 counter$count = 87382;
	#10 counter$count = 87383;
	#10 counter$count = 87384;
	#10 counter$count = 87385;
	#10 counter$count = 87386;
	#10 counter$count = 87387;
	#10 counter$count = 87388;
	#10 counter$count = 87389;
	#10 counter$count = 87390;
	#10 counter$count = 87391;
	#10 counter$count = 87392;
	#10 counter$count = 87393;
	#10 counter$count = 87394;
	#10 counter$count = 87395;
	#10 counter$count = 87396;
	#10 counter$count = 87397;
	#10 counter$count = 87398;
	#10 counter$count = 87399;
	#10 counter$count = 87400;
	#10 counter$count = 87401;
	#10 counter$count = 87402;
	#10 counter$count = 87403;
	#10 counter$count = 87404;
	#10 counter$count = 87405;
	#10 counter$count = 87406;
	#10 counter$count = 87407;
	#10 counter$count = 87408;
	#10 counter$count = 87409;
	#10 counter$count = 87410;
	#10 counter$count = 87411;
	#10 counter$count = 87412;
	#10 counter$count = 87413;
	#10 counter$count = 87414;
	#10 counter$count = 87415;
	#10 counter$count = 87416;
	#10 counter$count = 87417;
	#10 counter$count = 87418;
	#10 counter$count = 87419;
	#10 counter$count = 87420;
	#10 counter$count = 87421;
	#10 counter$count = 87422;
	#10 counter$count = 87423;
	#10 counter$count = 87424;
	#10 counter$count = 87425;
	#10 counter$count = 87426;
	#10 counter$count = 87427;
	#10 counter$count = 87428;
	#10 counter$count = 87429;
	#10 counter$count = 87430;
	#10 counter$count = 87431;
	#10 counter$count = 87432;
	#10 counter$count = 87433;
	#10 counter$count = 87434;
	#10 counter$count = 87435;
	#10 counter$count = 87436;
	#10 counter$count = 87437;
	#10 counter$count = 87438;
	#10 counter$count = 87439;
	#10 counter$count = 87440;
	#10 counter$count = 87441;
	#10 counter$count = 87442;
	#10 counter$count = 87443;
	#10 counter$count = 87444;
	#10 counter$count = 87445;
	#10 counter$count = 87446;
	#10 counter$count = 87447;
	#10 counter$count = 87448;
	#10 counter$count = 87449;
	#10 counter$count = 87450;
	#10 counter$count = 87451;
	#10 counter$count = 87452;
	#10 counter$count = 87453;
	#10 counter$count = 87454;
	#10 counter$count = 87455;
	#10 counter$count = 87456;
	#10 counter$count = 87457;
	#10 counter$count = 87458;
	#10 counter$count = 87459;
	#10 counter$count = 87460;
	#10 counter$count = 87461;
	#10 counter$count = 87462;
	#10 counter$count = 87463;
	#10 counter$count = 87464;
	#10 counter$count = 87465;
	#10 counter$count = 87466;
	#10 counter$count = 87467;
	#10 counter$count = 87468;
	#10 counter$count = 87469;
	#10 counter$count = 87470;
	#10 counter$count = 87471;
	#10 counter$count = 87472;
	#10 counter$count = 87473;
	#10 counter$count = 87474;
	#10 counter$count = 87475;
	#10 counter$count = 87476;
	#10 counter$count = 87477;
	#10 counter$count = 87478;
	#10 counter$count = 87479;
	#10 counter$count = 87480;
	#10 counter$count = 87481;
	#10 counter$count = 87482;
	#10 counter$count = 87483;
	#10 counter$count = 87484;
	#10 counter$count = 87485;
	#10 counter$count = 87486;
	#10 counter$count = 87487;
	#10 counter$count = 87488;
	#10 counter$count = 87489;
	#10 counter$count = 87490;
	#10 counter$count = 87491;
	#10 counter$count = 87492;
	#10 counter$count = 87493;
	#10 counter$count = 87494;
	#10 counter$count = 87495;
	#10 counter$count = 87496;
	#10 counter$count = 87497;
	#10 counter$count = 87498;
	#10 counter$count = 87499;
	#10 counter$count = 87500;
	#10 counter$count = 87501;
	#10 counter$count = 87502;
	#10 counter$count = 87503;
	#10 counter$count = 87504;
	#10 counter$count = 87505;
	#10 counter$count = 87506;
	#10 counter$count = 87507;
	#10 counter$count = 87508;
	#10 counter$count = 87509;
	#10 counter$count = 87510;
	#10 counter$count = 87511;
	#10 counter$count = 87512;
	#10 counter$count = 87513;
	#10 counter$count = 87514;
	#10 counter$count = 87515;
	#10 counter$count = 87516;
	#10 counter$count = 87517;
	#10 counter$count = 87518;
	#10 counter$count = 87519;
	#10 counter$count = 87520;
	#10 counter$count = 87521;
	#10 counter$count = 87522;
	#10 counter$count = 87523;
	#10 counter$count = 87524;
	#10 counter$count = 87525;
	#10 counter$count = 87526;
	#10 counter$count = 87527;
	#10 counter$count = 87528;
	#10 counter$count = 87529;
	#10 counter$count = 87530;
	#10 counter$count = 87531;
	#10 counter$count = 87532;
	#10 counter$count = 87533;
	#10 counter$count = 87534;
	#10 counter$count = 87535;
	#10 counter$count = 87536;
	#10 counter$count = 87537;
	#10 counter$count = 87538;
	#10 counter$count = 87539;
	#10 counter$count = 87540;
	#10 counter$count = 87541;
	#10 counter$count = 87542;
	#10 counter$count = 87543;
	#10 counter$count = 87544;
	#10 counter$count = 87545;
	#10 counter$count = 87546;
	#10 counter$count = 87547;
	#10 counter$count = 87548;
	#10 counter$count = 87549;
	#10 counter$count = 87550;
	#10 counter$count = 87551;
	#10 counter$count = 87552;
	#10 counter$count = 87553;
	#10 counter$count = 87554;
	#10 counter$count = 87555;
	#10 counter$count = 87556;
	#10 counter$count = 87557;
	#10 counter$count = 87558;
	#10 counter$count = 87559;
	#10 counter$count = 87560;
	#10 counter$count = 87561;
	#10 counter$count = 87562;
	#10 counter$count = 87563;
	#10 counter$count = 87564;
	#10 counter$count = 87565;
	#10 counter$count = 87566;
	#10 counter$count = 87567;
	#10 counter$count = 87568;
	#10 counter$count = 87569;
	#10 counter$count = 87570;
	#10 counter$count = 87571;
	#10 counter$count = 87572;
	#10 counter$count = 87573;
	#10 counter$count = 87574;
	#10 counter$count = 87575;
	#10 counter$count = 87576;
	#10 counter$count = 87577;
	#10 counter$count = 87578;
	#10 counter$count = 87579;
	#10 counter$count = 87580;
	#10 counter$count = 87581;
	#10 counter$count = 87582;
	#10 counter$count = 87583;
	#10 counter$count = 87584;
	#10 counter$count = 87585;
	#10 counter$count = 87586;
	#10 counter$count = 87587;
	#10 counter$count = 87588;
	#10 counter$count = 87589;
	#10 counter$count = 87590;
	#10 counter$count = 87591;
	#10 counter$count = 87592;
	#10 counter$count = 87593;
	#10 counter$count = 87594;
	#10 counter$count = 87595;
	#10 counter$count = 87596;
	#10 counter$count = 87597;
	#10 counter$count = 87598;
	#10 counter$count = 87599;
	#10 counter$count = 87600;
	#10 counter$count = 87601;
	#10 counter$count = 87602;
	#10 counter$count = 87603;
	#10 counter$count = 87604;
	#10 counter$count = 87605;
	#10 counter$count = 87606;
	#10 counter$count = 87607;
	#10 counter$count = 87608;
	#10 counter$count = 87609;
	#10 counter$count = 87610;
	#10 counter$count = 87611;
	#10 counter$count = 87612;
	#10 counter$count = 87613;
	#10 counter$count = 87614;
	#10 counter$count = 87615;
	#10 counter$count = 87616;
	#10 counter$count = 87617;
	#10 counter$count = 87618;
	#10 counter$count = 87619;
	#10 counter$count = 87620;
	#10 counter$count = 87621;
	#10 counter$count = 87622;
	#10 counter$count = 87623;
	#10 counter$count = 87624;
	#10 counter$count = 87625;
	#10 counter$count = 87626;
	#10 counter$count = 87627;
	#10 counter$count = 87628;
	#10 counter$count = 87629;
	#10 counter$count = 87630;
	#10 counter$count = 87631;
	#10 counter$count = 87632;
	#10 counter$count = 87633;
	#10 counter$count = 87634;
	#10 counter$count = 87635;
	#10 counter$count = 87636;
	#10 counter$count = 87637;
	#10 counter$count = 87638;
	#10 counter$count = 87639;
	#10 counter$count = 87640;
	#10 counter$count = 87641;
	#10 counter$count = 87642;
	#10 counter$count = 87643;
	#10 counter$count = 87644;
	#10 counter$count = 87645;
	#10 counter$count = 87646;
	#10 counter$count = 87647;
	#10 counter$count = 87648;
	#10 counter$count = 87649;
	#10 counter$count = 87650;
	#10 counter$count = 87651;
	#10 counter$count = 87652;
	#10 counter$count = 87653;
	#10 counter$count = 87654;
	#10 counter$count = 87655;
	#10 counter$count = 87656;
	#10 counter$count = 87657;
	#10 counter$count = 87658;
	#10 counter$count = 87659;
	#10 counter$count = 87660;
	#10 counter$count = 87661;
	#10 counter$count = 87662;
	#10 counter$count = 87663;
	#10 counter$count = 87664;
	#10 counter$count = 87665;
	#10 counter$count = 87666;
	#10 counter$count = 87667;
	#10 counter$count = 87668;
	#10 counter$count = 87669;
	#10 counter$count = 87670;
	#10 counter$count = 87671;
	#10 counter$count = 87672;
	#10 counter$count = 87673;
	#10 counter$count = 87674;
	#10 counter$count = 87675;
	#10 counter$count = 87676;
	#10 counter$count = 87677;
	#10 counter$count = 87678;
	#10 counter$count = 87679;
	#10 counter$count = 87680;
	#10 counter$count = 87681;
	#10 counter$count = 87682;
	#10 counter$count = 87683;
	#10 counter$count = 87684;
	#10 counter$count = 87685;
	#10 counter$count = 87686;
	#10 counter$count = 87687;
	#10 counter$count = 87688;
	#10 counter$count = 87689;
	#10 counter$count = 87690;
	#10 counter$count = 87691;
	#10 counter$count = 87692;
	#10 counter$count = 87693;
	#10 counter$count = 87694;
	#10 counter$count = 87695;
	#10 counter$count = 87696;
	#10 counter$count = 87697;
	#10 counter$count = 87698;
	#10 counter$count = 87699;
	#10 counter$count = 87700;
	#10 counter$count = 87701;
	#10 counter$count = 87702;
	#10 counter$count = 87703;
	#10 counter$count = 87704;
	#10 counter$count = 87705;
	#10 counter$count = 87706;
	#10 counter$count = 87707;
	#10 counter$count = 87708;
	#10 counter$count = 87709;
	#10 counter$count = 87710;
	#10 counter$count = 87711;
	#10 counter$count = 87712;
	#10 counter$count = 87713;
	#10 counter$count = 87714;
	#10 counter$count = 87715;
	#10 counter$count = 87716;
	#10 counter$count = 87717;
	#10 counter$count = 87718;
	#10 counter$count = 87719;
	#10 counter$count = 87720;
	#10 counter$count = 87721;
	#10 counter$count = 87722;
	#10 counter$count = 87723;
	#10 counter$count = 87724;
	#10 counter$count = 87725;
	#10 counter$count = 87726;
	#10 counter$count = 87727;
	#10 counter$count = 87728;
	#10 counter$count = 87729;
	#10 counter$count = 87730;
	#10 counter$count = 87731;
	#10 counter$count = 87732;
	#10 counter$count = 87733;
	#10 counter$count = 87734;
	#10 counter$count = 87735;
	#10 counter$count = 87736;
	#10 counter$count = 87737;
	#10 counter$count = 87738;
	#10 counter$count = 87739;
	#10 counter$count = 87740;
	#10 counter$count = 87741;
	#10 counter$count = 87742;
	#10 counter$count = 87743;
	#10 counter$count = 87744;
	#10 counter$count = 87745;
	#10 counter$count = 87746;
	#10 counter$count = 87747;
	#10 counter$count = 87748;
	#10 counter$count = 87749;
	#10 counter$count = 87750;
	#10 counter$count = 87751;
	#10 counter$count = 87752;
	#10 counter$count = 87753;
	#10 counter$count = 87754;
	#10 counter$count = 87755;
	#10 counter$count = 87756;
	#10 counter$count = 87757;
	#10 counter$count = 87758;
	#10 counter$count = 87759;
	#10 counter$count = 87760;
	#10 counter$count = 87761;
	#10 counter$count = 87762;
	#10 counter$count = 87763;
	#10 counter$count = 87764;
	#10 counter$count = 87765;
	#10 counter$count = 87766;
	#10 counter$count = 87767;
	#10 counter$count = 87768;
	#10 counter$count = 87769;
	#10 counter$count = 87770;
	#10 counter$count = 87771;
	#10 counter$count = 87772;
	#10 counter$count = 87773;
	#10 counter$count = 87774;
	#10 counter$count = 87775;
	#10 counter$count = 87776;
	#10 counter$count = 87777;
	#10 counter$count = 87778;
	#10 counter$count = 87779;
	#10 counter$count = 87780;
	#10 counter$count = 87781;
	#10 counter$count = 87782;
	#10 counter$count = 87783;
	#10 counter$count = 87784;
	#10 counter$count = 87785;
	#10 counter$count = 87786;
	#10 counter$count = 87787;
	#10 counter$count = 87788;
	#10 counter$count = 87789;
	#10 counter$count = 87790;
	#10 counter$count = 87791;
	#10 counter$count = 87792;
	#10 counter$count = 87793;
	#10 counter$count = 87794;
	#10 counter$count = 87795;
	#10 counter$count = 87796;
	#10 counter$count = 87797;
	#10 counter$count = 87798;
	#10 counter$count = 87799;
	#10 counter$count = 87800;
	#10 counter$count = 87801;
	#10 counter$count = 87802;
	#10 counter$count = 87803;
	#10 counter$count = 87804;
	#10 counter$count = 87805;
	#10 counter$count = 87806;
	#10 counter$count = 87807;
	#10 counter$count = 87808;
	#10 counter$count = 87809;
	#10 counter$count = 87810;
	#10 counter$count = 87811;
	#10 counter$count = 87812;
	#10 counter$count = 87813;
	#10 counter$count = 87814;
	#10 counter$count = 87815;
	#10 counter$count = 87816;
	#10 counter$count = 87817;
	#10 counter$count = 87818;
	#10 counter$count = 87819;
	#10 counter$count = 87820;
	#10 counter$count = 87821;
	#10 counter$count = 87822;
	#10 counter$count = 87823;
	#10 counter$count = 87824;
	#10 counter$count = 87825;
	#10 counter$count = 87826;
	#10 counter$count = 87827;
	#10 counter$count = 87828;
	#10 counter$count = 87829;
	#10 counter$count = 87830;
	#10 counter$count = 87831;
	#10 counter$count = 87832;
	#10 counter$count = 87833;
	#10 counter$count = 87834;
	#10 counter$count = 87835;
	#10 counter$count = 87836;
	#10 counter$count = 87837;
	#10 counter$count = 87838;
	#10 counter$count = 87839;
	#10 counter$count = 87840;
	#10 counter$count = 87841;
	#10 counter$count = 87842;
	#10 counter$count = 87843;
	#10 counter$count = 87844;
	#10 counter$count = 87845;
	#10 counter$count = 87846;
	#10 counter$count = 87847;
	#10 counter$count = 87848;
	#10 counter$count = 87849;
	#10 counter$count = 87850;
	#10 counter$count = 87851;
	#10 counter$count = 87852;
	#10 counter$count = 87853;
	#10 counter$count = 87854;
	#10 counter$count = 87855;
	#10 counter$count = 87856;
	#10 counter$count = 87857;
	#10 counter$count = 87858;
	#10 counter$count = 87859;
	#10 counter$count = 87860;
	#10 counter$count = 87861;
	#10 counter$count = 87862;
	#10 counter$count = 87863;
	#10 counter$count = 87864;
	#10 counter$count = 87865;
	#10 counter$count = 87866;
	#10 counter$count = 87867;
	#10 counter$count = 87868;
	#10 counter$count = 87869;
	#10 counter$count = 87870;
	#10 counter$count = 87871;
	#10 counter$count = 87872;
	#10 counter$count = 87873;
	#10 counter$count = 87874;
	#10 counter$count = 87875;
	#10 counter$count = 87876;
	#10 counter$count = 87877;
	#10 counter$count = 87878;
	#10 counter$count = 87879;
	#10 counter$count = 87880;
	#10 counter$count = 87881;
	#10 counter$count = 87882;
	#10 counter$count = 87883;
	#10 counter$count = 87884;
	#10 counter$count = 87885;
	#10 counter$count = 87886;
	#10 counter$count = 87887;
	#10 counter$count = 87888;
	#10 counter$count = 87889;
	#10 counter$count = 87890;
	#10 counter$count = 87891;
	#10 counter$count = 87892;
	#10 counter$count = 87893;
	#10 counter$count = 87894;
	#10 counter$count = 87895;
	#10 counter$count = 87896;
	#10 counter$count = 87897;
	#10 counter$count = 87898;
	#10 counter$count = 87899;
	#10 counter$count = 87900;
	#10 counter$count = 87901;
	#10 counter$count = 87902;
	#10 counter$count = 87903;
	#10 counter$count = 87904;
	#10 counter$count = 87905;
	#10 counter$count = 87906;
	#10 counter$count = 87907;
	#10 counter$count = 87908;
	#10 counter$count = 87909;
	#10 counter$count = 87910;
	#10 counter$count = 87911;
	#10 counter$count = 87912;
	#10 counter$count = 87913;
	#10 counter$count = 87914;
	#10 counter$count = 87915;
	#10 counter$count = 87916;
	#10 counter$count = 87917;
	#10 counter$count = 87918;
	#10 counter$count = 87919;
	#10 counter$count = 87920;
	#10 counter$count = 87921;
	#10 counter$count = 87922;
	#10 counter$count = 87923;
	#10 counter$count = 87924;
	#10 counter$count = 87925;
	#10 counter$count = 87926;
	#10 counter$count = 87927;
	#10 counter$count = 87928;
	#10 counter$count = 87929;
	#10 counter$count = 87930;
	#10 counter$count = 87931;
	#10 counter$count = 87932;
	#10 counter$count = 87933;
	#10 counter$count = 87934;
	#10 counter$count = 87935;
	#10 counter$count = 87936;
	#10 counter$count = 87937;
	#10 counter$count = 87938;
	#10 counter$count = 87939;
	#10 counter$count = 87940;
	#10 counter$count = 87941;
	#10 counter$count = 87942;
	#10 counter$count = 87943;
	#10 counter$count = 87944;
	#10 counter$count = 87945;
	#10 counter$count = 87946;
	#10 counter$count = 87947;
	#10 counter$count = 87948;
	#10 counter$count = 87949;
	#10 counter$count = 87950;
	#10 counter$count = 87951;
	#10 counter$count = 87952;
	#10 counter$count = 87953;
	#10 counter$count = 87954;
	#10 counter$count = 87955;
	#10 counter$count = 87956;
	#10 counter$count = 87957;
	#10 counter$count = 87958;
	#10 counter$count = 87959;
	#10 counter$count = 87960;
	#10 counter$count = 87961;
	#10 counter$count = 87962;
	#10 counter$count = 87963;
	#10 counter$count = 87964;
	#10 counter$count = 87965;
	#10 counter$count = 87966;
	#10 counter$count = 87967;
	#10 counter$count = 87968;
	#10 counter$count = 87969;
	#10 counter$count = 87970;
	#10 counter$count = 87971;
	#10 counter$count = 87972;
	#10 counter$count = 87973;
	#10 counter$count = 87974;
	#10 counter$count = 87975;
	#10 counter$count = 87976;
	#10 counter$count = 87977;
	#10 counter$count = 87978;
	#10 counter$count = 87979;
	#10 counter$count = 87980;
	#10 counter$count = 87981;
	#10 counter$count = 87982;
	#10 counter$count = 87983;
	#10 counter$count = 87984;
	#10 counter$count = 87985;
	#10 counter$count = 87986;
	#10 counter$count = 87987;
	#10 counter$count = 87988;
	#10 counter$count = 87989;
	#10 counter$count = 87990;
	#10 counter$count = 87991;
	#10 counter$count = 87992;
	#10 counter$count = 87993;
	#10 counter$count = 87994;
	#10 counter$count = 87995;
	#10 counter$count = 87996;
	#10 counter$count = 87997;
	#10 counter$count = 87998;
	#10 counter$count = 87999;
	#10 counter$count = 88000;
	#10 counter$count = 88001;
	#10 counter$count = 88002;
	#10 counter$count = 88003;
	#10 counter$count = 88004;
	#10 counter$count = 88005;
	#10 counter$count = 88006;
	#10 counter$count = 88007;
	#10 counter$count = 88008;
	#10 counter$count = 88009;
	#10 counter$count = 88010;
	#10 counter$count = 88011;
	#10 counter$count = 88012;
	#10 counter$count = 88013;
	#10 counter$count = 88014;
	#10 counter$count = 88015;
	#10 counter$count = 88016;
	#10 counter$count = 88017;
	#10 counter$count = 88018;
	#10 counter$count = 88019;
	#10 counter$count = 88020;
	#10 counter$count = 88021;
	#10 counter$count = 88022;
	#10 counter$count = 88023;
	#10 counter$count = 88024;
	#10 counter$count = 88025;
	#10 counter$count = 88026;
	#10 counter$count = 88027;
	#10 counter$count = 88028;
	#10 counter$count = 88029;
	#10 counter$count = 88030;
	#10 counter$count = 88031;
	#10 counter$count = 88032;
	#10 counter$count = 88033;
	#10 counter$count = 88034;
	#10 counter$count = 88035;
	#10 counter$count = 88036;
	#10 counter$count = 88037;
	#10 counter$count = 88038;
	#10 counter$count = 88039;
	#10 counter$count = 88040;
	#10 counter$count = 88041;
	#10 counter$count = 88042;
	#10 counter$count = 88043;
	#10 counter$count = 88044;
	#10 counter$count = 88045;
	#10 counter$count = 88046;
	#10 counter$count = 88047;
	#10 counter$count = 88048;
	#10 counter$count = 88049;
	#10 counter$count = 88050;
	#10 counter$count = 88051;
	#10 counter$count = 88052;
	#10 counter$count = 88053;
	#10 counter$count = 88054;
	#10 counter$count = 88055;
	#10 counter$count = 88056;
	#10 counter$count = 88057;
	#10 counter$count = 88058;
	#10 counter$count = 88059;
	#10 counter$count = 88060;
	#10 counter$count = 88061;
	#10 counter$count = 88062;
	#10 counter$count = 88063;
	#10 counter$count = 88064;
	#10 counter$count = 88065;
	#10 counter$count = 88066;
	#10 counter$count = 88067;
	#10 counter$count = 88068;
	#10 counter$count = 88069;
	#10 counter$count = 88070;
	#10 counter$count = 88071;
	#10 counter$count = 88072;
	#10 counter$count = 88073;
	#10 counter$count = 88074;
	#10 counter$count = 88075;
	#10 counter$count = 88076;
	#10 counter$count = 88077;
	#10 counter$count = 88078;
	#10 counter$count = 88079;
	#10 counter$count = 88080;
	#10 counter$count = 88081;
	#10 counter$count = 88082;
	#10 counter$count = 88083;
	#10 counter$count = 88084;
	#10 counter$count = 88085;
	#10 counter$count = 88086;
	#10 counter$count = 88087;
	#10 counter$count = 88088;
	#10 counter$count = 88089;
	#10 counter$count = 88090;
	#10 counter$count = 88091;
	#10 counter$count = 88092;
	#10 counter$count = 88093;
	#10 counter$count = 88094;
	#10 counter$count = 88095;
	#10 counter$count = 88096;
	#10 counter$count = 88097;
	#10 counter$count = 88098;
	#10 counter$count = 88099;
	#10 counter$count = 88100;
	#10 counter$count = 88101;
	#10 counter$count = 88102;
	#10 counter$count = 88103;
	#10 counter$count = 88104;
	#10 counter$count = 88105;
	#10 counter$count = 88106;
	#10 counter$count = 88107;
	#10 counter$count = 88108;
	#10 counter$count = 88109;
	#10 counter$count = 88110;
	#10 counter$count = 88111;
	#10 counter$count = 88112;
	#10 counter$count = 88113;
	#10 counter$count = 88114;
	#10 counter$count = 88115;
	#10 counter$count = 88116;
	#10 counter$count = 88117;
	#10 counter$count = 88118;
	#10 counter$count = 88119;
	#10 counter$count = 88120;
	#10 counter$count = 88121;
	#10 counter$count = 88122;
	#10 counter$count = 88123;
	#10 counter$count = 88124;
	#10 counter$count = 88125;
	#10 counter$count = 88126;
	#10 counter$count = 88127;
	#10 counter$count = 88128;
	#10 counter$count = 88129;
	#10 counter$count = 88130;
	#10 counter$count = 88131;
	#10 counter$count = 88132;
	#10 counter$count = 88133;
	#10 counter$count = 88134;
	#10 counter$count = 88135;
	#10 counter$count = 88136;
	#10 counter$count = 88137;
	#10 counter$count = 88138;
	#10 counter$count = 88139;
	#10 counter$count = 88140;
	#10 counter$count = 88141;
	#10 counter$count = 88142;
	#10 counter$count = 88143;
	#10 counter$count = 88144;
	#10 counter$count = 88145;
	#10 counter$count = 88146;
	#10 counter$count = 88147;
	#10 counter$count = 88148;
	#10 counter$count = 88149;
	#10 counter$count = 88150;
	#10 counter$count = 88151;
	#10 counter$count = 88152;
	#10 counter$count = 88153;
	#10 counter$count = 88154;
	#10 counter$count = 88155;
	#10 counter$count = 88156;
	#10 counter$count = 88157;
	#10 counter$count = 88158;
	#10 counter$count = 88159;
	#10 counter$count = 88160;
	#10 counter$count = 88161;
	#10 counter$count = 88162;
	#10 counter$count = 88163;
	#10 counter$count = 88164;
	#10 counter$count = 88165;
	#10 counter$count = 88166;
	#10 counter$count = 88167;
	#10 counter$count = 88168;
	#10 counter$count = 88169;
	#10 counter$count = 88170;
	#10 counter$count = 88171;
	#10 counter$count = 88172;
	#10 counter$count = 88173;
	#10 counter$count = 88174;
	#10 counter$count = 88175;
	#10 counter$count = 88176;
	#10 counter$count = 88177;
	#10 counter$count = 88178;
	#10 counter$count = 88179;
	#10 counter$count = 88180;
	#10 counter$count = 88181;
	#10 counter$count = 88182;
	#10 counter$count = 88183;
	#10 counter$count = 88184;
	#10 counter$count = 88185;
	#10 counter$count = 88186;
	#10 counter$count = 88187;
	#10 counter$count = 88188;
	#10 counter$count = 88189;
	#10 counter$count = 88190;
	#10 counter$count = 88191;
	#10 counter$count = 88192;
	#10 counter$count = 88193;
	#10 counter$count = 88194;
	#10 counter$count = 88195;
	#10 counter$count = 88196;
	#10 counter$count = 88197;
	#10 counter$count = 88198;
	#10 counter$count = 88199;
	#10 counter$count = 88200;
	#10 counter$count = 88201;
	#10 counter$count = 88202;
	#10 counter$count = 88203;
	#10 counter$count = 88204;
	#10 counter$count = 88205;
	#10 counter$count = 88206;
	#10 counter$count = 88207;
	#10 counter$count = 88208;
	#10 counter$count = 88209;
	#10 counter$count = 88210;
	#10 counter$count = 88211;
	#10 counter$count = 88212;
	#10 counter$count = 88213;
	#10 counter$count = 88214;
	#10 counter$count = 88215;
	#10 counter$count = 88216;
	#10 counter$count = 88217;
	#10 counter$count = 88218;
	#10 counter$count = 88219;
	#10 counter$count = 88220;
	#10 counter$count = 88221;
	#10 counter$count = 88222;
	#10 counter$count = 88223;
	#10 counter$count = 88224;
	#10 counter$count = 88225;
	#10 counter$count = 88226;
	#10 counter$count = 88227;
	#10 counter$count = 88228;
	#10 counter$count = 88229;
	#10 counter$count = 88230;
	#10 counter$count = 88231;
	#10 counter$count = 88232;
	#10 counter$count = 88233;
	#10 counter$count = 88234;
	#10 counter$count = 88235;
	#10 counter$count = 88236;
	#10 counter$count = 88237;
	#10 counter$count = 88238;
	#10 counter$count = 88239;
	#10 counter$count = 88240;
	#10 counter$count = 88241;
	#10 counter$count = 88242;
	#10 counter$count = 88243;
	#10 counter$count = 88244;
	#10 counter$count = 88245;
	#10 counter$count = 88246;
	#10 counter$count = 88247;
	#10 counter$count = 88248;
	#10 counter$count = 88249;
	#10 counter$count = 88250;
	#10 counter$count = 88251;
	#10 counter$count = 88252;
	#10 counter$count = 88253;
	#10 counter$count = 88254;
	#10 counter$count = 88255;
	#10 counter$count = 88256;
	#10 counter$count = 88257;
	#10 counter$count = 88258;
	#10 counter$count = 88259;
	#10 counter$count = 88260;
	#10 counter$count = 88261;
	#10 counter$count = 88262;
	#10 counter$count = 88263;
	#10 counter$count = 88264;
	#10 counter$count = 88265;
	#10 counter$count = 88266;
	#10 counter$count = 88267;
	#10 counter$count = 88268;
	#10 counter$count = 88269;
	#10 counter$count = 88270;
	#10 counter$count = 88271;
	#10 counter$count = 88272;
	#10 counter$count = 88273;
	#10 counter$count = 88274;
	#10 counter$count = 88275;
	#10 counter$count = 88276;
	#10 counter$count = 88277;
	#10 counter$count = 88278;
	#10 counter$count = 88279;
	#10 counter$count = 88280;
	#10 counter$count = 88281;
	#10 counter$count = 88282;
	#10 counter$count = 88283;
	#10 counter$count = 88284;
	#10 counter$count = 88285;
	#10 counter$count = 88286;
	#10 counter$count = 88287;
	#10 counter$count = 88288;
	#10 counter$count = 88289;
	#10 counter$count = 88290;
	#10 counter$count = 88291;
	#10 counter$count = 88292;
	#10 counter$count = 88293;
	#10 counter$count = 88294;
	#10 counter$count = 88295;
	#10 counter$count = 88296;
	#10 counter$count = 88297;
	#10 counter$count = 88298;
	#10 counter$count = 88299;
	#10 counter$count = 88300;
	#10 counter$count = 88301;
	#10 counter$count = 88302;
	#10 counter$count = 88303;
	#10 counter$count = 88304;
	#10 counter$count = 88305;
	#10 counter$count = 88306;
	#10 counter$count = 88307;
	#10 counter$count = 88308;
	#10 counter$count = 88309;
	#10 counter$count = 88310;
	#10 counter$count = 88311;
	#10 counter$count = 88312;
	#10 counter$count = 88313;
	#10 counter$count = 88314;
	#10 counter$count = 88315;
	#10 counter$count = 88316;
	#10 counter$count = 88317;
	#10 counter$count = 88318;
	#10 counter$count = 88319;
	#10 counter$count = 88320;
	#10 counter$count = 88321;
	#10 counter$count = 88322;
	#10 counter$count = 88323;
	#10 counter$count = 88324;
	#10 counter$count = 88325;
	#10 counter$count = 88326;
	#10 counter$count = 88327;
	#10 counter$count = 88328;
	#10 counter$count = 88329;
	#10 counter$count = 88330;
	#10 counter$count = 88331;
	#10 counter$count = 88332;
	#10 counter$count = 88333;
	#10 counter$count = 88334;
	#10 counter$count = 88335;
	#10 counter$count = 88336;
	#10 counter$count = 88337;
	#10 counter$count = 88338;
	#10 counter$count = 88339;
	#10 counter$count = 88340;
	#10 counter$count = 88341;
	#10 counter$count = 88342;
	#10 counter$count = 88343;
	#10 counter$count = 88344;
	#10 counter$count = 88345;
	#10 counter$count = 88346;
	#10 counter$count = 88347;
	#10 counter$count = 88348;
	#10 counter$count = 88349;
	#10 counter$count = 88350;
	#10 counter$count = 88351;
	#10 counter$count = 88352;
	#10 counter$count = 88353;
	#10 counter$count = 88354;
	#10 counter$count = 88355;
	#10 counter$count = 88356;
	#10 counter$count = 88357;
	#10 counter$count = 88358;
	#10 counter$count = 88359;
	#10 counter$count = 88360;
	#10 counter$count = 88361;
	#10 counter$count = 88362;
	#10 counter$count = 88363;
	#10 counter$count = 88364;
	#10 counter$count = 88365;
	#10 counter$count = 88366;
	#10 counter$count = 88367;
	#10 counter$count = 88368;
	#10 counter$count = 88369;
	#10 counter$count = 88370;
	#10 counter$count = 88371;
	#10 counter$count = 88372;
	#10 counter$count = 88373;
	#10 counter$count = 88374;
	#10 counter$count = 88375;
	#10 counter$count = 88376;
	#10 counter$count = 88377;
	#10 counter$count = 88378;
	#10 counter$count = 88379;
	#10 counter$count = 88380;
	#10 counter$count = 88381;
	#10 counter$count = 88382;
	#10 counter$count = 88383;
	#10 counter$count = 88384;
	#10 counter$count = 88385;
	#10 counter$count = 88386;
	#10 counter$count = 88387;
	#10 counter$count = 88388;
	#10 counter$count = 88389;
	#10 counter$count = 88390;
	#10 counter$count = 88391;
	#10 counter$count = 88392;
	#10 counter$count = 88393;
	#10 counter$count = 88394;
	#10 counter$count = 88395;
	#10 counter$count = 88396;
	#10 counter$count = 88397;
	#10 counter$count = 88398;
	#10 counter$count = 88399;
	#10 counter$count = 88400;
	#10 counter$count = 88401;
	#10 counter$count = 88402;
	#10 counter$count = 88403;
	#10 counter$count = 88404;
	#10 counter$count = 88405;
	#10 counter$count = 88406;
	#10 counter$count = 88407;
	#10 counter$count = 88408;
	#10 counter$count = 88409;
	#10 counter$count = 88410;
	#10 counter$count = 88411;
	#10 counter$count = 88412;
	#10 counter$count = 88413;
	#10 counter$count = 88414;
	#10 counter$count = 88415;
	#10 counter$count = 88416;
	#10 counter$count = 88417;
	#10 counter$count = 88418;
	#10 counter$count = 88419;
	#10 counter$count = 88420;
	#10 counter$count = 88421;
	#10 counter$count = 88422;
	#10 counter$count = 88423;
	#10 counter$count = 88424;
	#10 counter$count = 88425;
	#10 counter$count = 88426;
	#10 counter$count = 88427;
	#10 counter$count = 88428;
	#10 counter$count = 88429;
	#10 counter$count = 88430;
	#10 counter$count = 88431;
	#10 counter$count = 88432;
	#10 counter$count = 88433;
	#10 counter$count = 88434;
	#10 counter$count = 88435;
	#10 counter$count = 88436;
	#10 counter$count = 88437;
	#10 counter$count = 88438;
	#10 counter$count = 88439;
	#10 counter$count = 88440;
	#10 counter$count = 88441;
	#10 counter$count = 88442;
	#10 counter$count = 88443;
	#10 counter$count = 88444;
	#10 counter$count = 88445;
	#10 counter$count = 88446;
	#10 counter$count = 88447;
	#10 counter$count = 88448;
	#10 counter$count = 88449;
	#10 counter$count = 88450;
	#10 counter$count = 88451;
	#10 counter$count = 88452;
	#10 counter$count = 88453;
	#10 counter$count = 88454;
	#10 counter$count = 88455;
	#10 counter$count = 88456;
	#10 counter$count = 88457;
	#10 counter$count = 88458;
	#10 counter$count = 88459;
	#10 counter$count = 88460;
	#10 counter$count = 88461;
	#10 counter$count = 88462;
	#10 counter$count = 88463;
	#10 counter$count = 88464;
	#10 counter$count = 88465;
	#10 counter$count = 88466;
	#10 counter$count = 88467;
	#10 counter$count = 88468;
	#10 counter$count = 88469;
	#10 counter$count = 88470;
	#10 counter$count = 88471;
	#10 counter$count = 88472;
	#10 counter$count = 88473;
	#10 counter$count = 88474;
	#10 counter$count = 88475;
	#10 counter$count = 88476;
	#10 counter$count = 88477;
	#10 counter$count = 88478;
	#10 counter$count = 88479;
	#10 counter$count = 88480;
	#10 counter$count = 88481;
	#10 counter$count = 88482;
	#10 counter$count = 88483;
	#10 counter$count = 88484;
	#10 counter$count = 88485;
	#10 counter$count = 88486;
	#10 counter$count = 88487;
	#10 counter$count = 88488;
	#10 counter$count = 88489;
	#10 counter$count = 88490;
	#10 counter$count = 88491;
	#10 counter$count = 88492;
	#10 counter$count = 88493;
	#10 counter$count = 88494;
	#10 counter$count = 88495;
	#10 counter$count = 88496;
	#10 counter$count = 88497;
	#10 counter$count = 88498;
	#10 counter$count = 88499;
	#10 counter$count = 88500;
	#10 counter$count = 88501;
	#10 counter$count = 88502;
	#10 counter$count = 88503;
	#10 counter$count = 88504;
	#10 counter$count = 88505;
	#10 counter$count = 88506;
	#10 counter$count = 88507;
	#10 counter$count = 88508;
	#10 counter$count = 88509;
	#10 counter$count = 88510;
	#10 counter$count = 88511;
	#10 counter$count = 88512;
	#10 counter$count = 88513;
	#10 counter$count = 88514;
	#10 counter$count = 88515;
	#10 counter$count = 88516;
	#10 counter$count = 88517;
	#10 counter$count = 88518;
	#10 counter$count = 88519;
	#10 counter$count = 88520;
	#10 counter$count = 88521;
	#10 counter$count = 88522;
	#10 counter$count = 88523;
	#10 counter$count = 88524;
	#10 counter$count = 88525;
	#10 counter$count = 88526;
	#10 counter$count = 88527;
	#10 counter$count = 88528;
	#10 counter$count = 88529;
	#10 counter$count = 88530;
	#10 counter$count = 88531;
	#10 counter$count = 88532;
	#10 counter$count = 88533;
	#10 counter$count = 88534;
	#10 counter$count = 88535;
	#10 counter$count = 88536;
	#10 counter$count = 88537;
	#10 counter$count = 88538;
	#10 counter$count = 88539;
	#10 counter$count = 88540;
	#10 counter$count = 88541;
	#10 counter$count = 88542;
	#10 counter$count = 88543;
	#10 counter$count = 88544;
	#10 counter$count = 88545;
	#10 counter$count = 88546;
	#10 counter$count = 88547;
	#10 counter$count = 88548;
	#10 counter$count = 88549;
	#10 counter$count = 88550;
	#10 counter$count = 88551;
	#10 counter$count = 88552;
	#10 counter$count = 88553;
	#10 counter$count = 88554;
	#10 counter$count = 88555;
	#10 counter$count = 88556;
	#10 counter$count = 88557;
	#10 counter$count = 88558;
	#10 counter$count = 88559;
	#10 counter$count = 88560;
	#10 counter$count = 88561;
	#10 counter$count = 88562;
	#10 counter$count = 88563;
	#10 counter$count = 88564;
	#10 counter$count = 88565;
	#10 counter$count = 88566;
	#10 counter$count = 88567;
	#10 counter$count = 88568;
	#10 counter$count = 88569;
	#10 counter$count = 88570;
	#10 counter$count = 88571;
	#10 counter$count = 88572;
	#10 counter$count = 88573;
	#10 counter$count = 88574;
	#10 counter$count = 88575;
	#10 counter$count = 88576;
	#10 counter$count = 88577;
	#10 counter$count = 88578;
	#10 counter$count = 88579;
	#10 counter$count = 88580;
	#10 counter$count = 88581;
	#10 counter$count = 88582;
	#10 counter$count = 88583;
	#10 counter$count = 88584;
	#10 counter$count = 88585;
	#10 counter$count = 88586;
	#10 counter$count = 88587;
	#10 counter$count = 88588;
	#10 counter$count = 88589;
	#10 counter$count = 88590;
	#10 counter$count = 88591;
	#10 counter$count = 88592;
	#10 counter$count = 88593;
	#10 counter$count = 88594;
	#10 counter$count = 88595;
	#10 counter$count = 88596;
	#10 counter$count = 88597;
	#10 counter$count = 88598;
	#10 counter$count = 88599;
	#10 counter$count = 88600;
	#10 counter$count = 88601;
	#10 counter$count = 88602;
	#10 counter$count = 88603;
	#10 counter$count = 88604;
	#10 counter$count = 88605;
	#10 counter$count = 88606;
	#10 counter$count = 88607;
	#10 counter$count = 88608;
	#10 counter$count = 88609;
	#10 counter$count = 88610;
	#10 counter$count = 88611;
	#10 counter$count = 88612;
	#10 counter$count = 88613;
	#10 counter$count = 88614;
	#10 counter$count = 88615;
	#10 counter$count = 88616;
	#10 counter$count = 88617;
	#10 counter$count = 88618;
	#10 counter$count = 88619;
	#10 counter$count = 88620;
	#10 counter$count = 88621;
	#10 counter$count = 88622;
	#10 counter$count = 88623;
	#10 counter$count = 88624;
	#10 counter$count = 88625;
	#10 counter$count = 88626;
	#10 counter$count = 88627;
	#10 counter$count = 88628;
	#10 counter$count = 88629;
	#10 counter$count = 88630;
	#10 counter$count = 88631;
	#10 counter$count = 88632;
	#10 counter$count = 88633;
	#10 counter$count = 88634;
	#10 counter$count = 88635;
	#10 counter$count = 88636;
	#10 counter$count = 88637;
	#10 counter$count = 88638;
	#10 counter$count = 88639;
	#10 counter$count = 88640;
	#10 counter$count = 88641;
	#10 counter$count = 88642;
	#10 counter$count = 88643;
	#10 counter$count = 88644;
	#10 counter$count = 88645;
	#10 counter$count = 88646;
	#10 counter$count = 88647;
	#10 counter$count = 88648;
	#10 counter$count = 88649;
	#10 counter$count = 88650;
	#10 counter$count = 88651;
	#10 counter$count = 88652;
	#10 counter$count = 88653;
	#10 counter$count = 88654;
	#10 counter$count = 88655;
	#10 counter$count = 88656;
	#10 counter$count = 88657;
	#10 counter$count = 88658;
	#10 counter$count = 88659;
	#10 counter$count = 88660;
	#10 counter$count = 88661;
	#10 counter$count = 88662;
	#10 counter$count = 88663;
	#10 counter$count = 88664;
	#10 counter$count = 88665;
	#10 counter$count = 88666;
	#10 counter$count = 88667;
	#10 counter$count = 88668;
	#10 counter$count = 88669;
	#10 counter$count = 88670;
	#10 counter$count = 88671;
	#10 counter$count = 88672;
	#10 counter$count = 88673;
	#10 counter$count = 88674;
	#10 counter$count = 88675;
	#10 counter$count = 88676;
	#10 counter$count = 88677;
	#10 counter$count = 88678;
	#10 counter$count = 88679;
	#10 counter$count = 88680;
	#10 counter$count = 88681;
	#10 counter$count = 88682;
	#10 counter$count = 88683;
	#10 counter$count = 88684;
	#10 counter$count = 88685;
	#10 counter$count = 88686;
	#10 counter$count = 88687;
	#10 counter$count = 88688;
	#10 counter$count = 88689;
	#10 counter$count = 88690;
	#10 counter$count = 88691;
	#10 counter$count = 88692;
	#10 counter$count = 88693;
	#10 counter$count = 88694;
	#10 counter$count = 88695;
	#10 counter$count = 88696;
	#10 counter$count = 88697;
	#10 counter$count = 88698;
	#10 counter$count = 88699;
	#10 counter$count = 88700;
	#10 counter$count = 88701;
	#10 counter$count = 88702;
	#10 counter$count = 88703;
	#10 counter$count = 88704;
	#10 counter$count = 88705;
	#10 counter$count = 88706;
	#10 counter$count = 88707;
	#10 counter$count = 88708;
	#10 counter$count = 88709;
	#10 counter$count = 88710;
	#10 counter$count = 88711;
	#10 counter$count = 88712;
	#10 counter$count = 88713;
	#10 counter$count = 88714;
	#10 counter$count = 88715;
	#10 counter$count = 88716;
	#10 counter$count = 88717;
	#10 counter$count = 88718;
	#10 counter$count = 88719;
	#10 counter$count = 88720;
	#10 counter$count = 88721;
	#10 counter$count = 88722;
	#10 counter$count = 88723;
	#10 counter$count = 88724;
	#10 counter$count = 88725;
	#10 counter$count = 88726;
	#10 counter$count = 88727;
	#10 counter$count = 88728;
	#10 counter$count = 88729;
	#10 counter$count = 88730;
	#10 counter$count = 88731;
	#10 counter$count = 88732;
	#10 counter$count = 88733;
	#10 counter$count = 88734;
	#10 counter$count = 88735;
	#10 counter$count = 88736;
	#10 counter$count = 88737;
	#10 counter$count = 88738;
	#10 counter$count = 88739;
	#10 counter$count = 88740;
	#10 counter$count = 88741;
	#10 counter$count = 88742;
	#10 counter$count = 88743;
	#10 counter$count = 88744;
	#10 counter$count = 88745;
	#10 counter$count = 88746;
	#10 counter$count = 88747;
	#10 counter$count = 88748;
	#10 counter$count = 88749;
	#10 counter$count = 88750;
	#10 counter$count = 88751;
	#10 counter$count = 88752;
	#10 counter$count = 88753;
	#10 counter$count = 88754;
	#10 counter$count = 88755;
	#10 counter$count = 88756;
	#10 counter$count = 88757;
	#10 counter$count = 88758;
	#10 counter$count = 88759;
	#10 counter$count = 88760;
	#10 counter$count = 88761;
	#10 counter$count = 88762;
	#10 counter$count = 88763;
	#10 counter$count = 88764;
	#10 counter$count = 88765;
	#10 counter$count = 88766;
	#10 counter$count = 88767;
	#10 counter$count = 88768;
	#10 counter$count = 88769;
	#10 counter$count = 88770;
	#10 counter$count = 88771;
	#10 counter$count = 88772;
	#10 counter$count = 88773;
	#10 counter$count = 88774;
	#10 counter$count = 88775;
	#10 counter$count = 88776;
	#10 counter$count = 88777;
	#10 counter$count = 88778;
	#10 counter$count = 88779;
	#10 counter$count = 88780;
	#10 counter$count = 88781;
	#10 counter$count = 88782;
	#10 counter$count = 88783;
	#10 counter$count = 88784;
	#10 counter$count = 88785;
	#10 counter$count = 88786;
	#10 counter$count = 88787;
	#10 counter$count = 88788;
	#10 counter$count = 88789;
	#10 counter$count = 88790;
	#10 counter$count = 88791;
	#10 counter$count = 88792;
	#10 counter$count = 88793;
	#10 counter$count = 88794;
	#10 counter$count = 88795;
	#10 counter$count = 88796;
	#10 counter$count = 88797;
	#10 counter$count = 88798;
	#10 counter$count = 88799;
	#10 counter$count = 88800;
	#10 counter$count = 88801;
	#10 counter$count = 88802;
	#10 counter$count = 88803;
	#10 counter$count = 88804;
	#10 counter$count = 88805;
	#10 counter$count = 88806;
	#10 counter$count = 88807;
	#10 counter$count = 88808;
	#10 counter$count = 88809;
	#10 counter$count = 88810;
	#10 counter$count = 88811;
	#10 counter$count = 88812;
	#10 counter$count = 88813;
	#10 counter$count = 88814;
	#10 counter$count = 88815;
	#10 counter$count = 88816;
	#10 counter$count = 88817;
	#10 counter$count = 88818;
	#10 counter$count = 88819;
	#10 counter$count = 88820;
	#10 counter$count = 88821;
	#10 counter$count = 88822;
	#10 counter$count = 88823;
	#10 counter$count = 88824;
	#10 counter$count = 88825;
	#10 counter$count = 88826;
	#10 counter$count = 88827;
	#10 counter$count = 88828;
	#10 counter$count = 88829;
	#10 counter$count = 88830;
	#10 counter$count = 88831;
	#10 counter$count = 88832;
	#10 counter$count = 88833;
	#10 counter$count = 88834;
	#10 counter$count = 88835;
	#10 counter$count = 88836;
	#10 counter$count = 88837;
	#10 counter$count = 88838;
	#10 counter$count = 88839;
	#10 counter$count = 88840;
	#10 counter$count = 88841;
	#10 counter$count = 88842;
	#10 counter$count = 88843;
	#10 counter$count = 88844;
	#10 counter$count = 88845;
	#10 counter$count = 88846;
	#10 counter$count = 88847;
	#10 counter$count = 88848;
	#10 counter$count = 88849;
	#10 counter$count = 88850;
	#10 counter$count = 88851;
	#10 counter$count = 88852;
	#10 counter$count = 88853;
	#10 counter$count = 88854;
	#10 counter$count = 88855;
	#10 counter$count = 88856;
	#10 counter$count = 88857;
	#10 counter$count = 88858;
	#10 counter$count = 88859;
	#10 counter$count = 88860;
	#10 counter$count = 88861;
	#10 counter$count = 88862;
	#10 counter$count = 88863;
	#10 counter$count = 88864;
	#10 counter$count = 88865;
	#10 counter$count = 88866;
	#10 counter$count = 88867;
	#10 counter$count = 88868;
	#10 counter$count = 88869;
	#10 counter$count = 88870;
	#10 counter$count = 88871;
	#10 counter$count = 88872;
	#10 counter$count = 88873;
	#10 counter$count = 88874;
	#10 counter$count = 88875;
	#10 counter$count = 88876;
	#10 counter$count = 88877;
	#10 counter$count = 88878;
	#10 counter$count = 88879;
	#10 counter$count = 88880;
	#10 counter$count = 88881;
	#10 counter$count = 88882;
	#10 counter$count = 88883;
	#10 counter$count = 88884;
	#10 counter$count = 88885;
	#10 counter$count = 88886;
	#10 counter$count = 88887;
	#10 counter$count = 88888;
	#10 counter$count = 88889;
	#10 counter$count = 88890;
	#10 counter$count = 88891;
	#10 counter$count = 88892;
	#10 counter$count = 88893;
	#10 counter$count = 88894;
	#10 counter$count = 88895;
	#10 counter$count = 88896;
	#10 counter$count = 88897;
	#10 counter$count = 88898;
	#10 counter$count = 88899;
	#10 counter$count = 88900;
	#10 counter$count = 88901;
	#10 counter$count = 88902;
	#10 counter$count = 88903;
	#10 counter$count = 88904;
	#10 counter$count = 88905;
	#10 counter$count = 88906;
	#10 counter$count = 88907;
	#10 counter$count = 88908;
	#10 counter$count = 88909;
	#10 counter$count = 88910;
	#10 counter$count = 88911;
	#10 counter$count = 88912;
	#10 counter$count = 88913;
	#10 counter$count = 88914;
	#10 counter$count = 88915;
	#10 counter$count = 88916;
	#10 counter$count = 88917;
	#10 counter$count = 88918;
	#10 counter$count = 88919;
	#10 counter$count = 88920;
	#10 counter$count = 88921;
	#10 counter$count = 88922;
	#10 counter$count = 88923;
	#10 counter$count = 88924;
	#10 counter$count = 88925;
	#10 counter$count = 88926;
	#10 counter$count = 88927;
	#10 counter$count = 88928;
	#10 counter$count = 88929;
	#10 counter$count = 88930;
	#10 counter$count = 88931;
	#10 counter$count = 88932;
	#10 counter$count = 88933;
	#10 counter$count = 88934;
	#10 counter$count = 88935;
	#10 counter$count = 88936;
	#10 counter$count = 88937;
	#10 counter$count = 88938;
	#10 counter$count = 88939;
	#10 counter$count = 88940;
	#10 counter$count = 88941;
	#10 counter$count = 88942;
	#10 counter$count = 88943;
	#10 counter$count = 88944;
	#10 counter$count = 88945;
	#10 counter$count = 88946;
	#10 counter$count = 88947;
	#10 counter$count = 88948;
	#10 counter$count = 88949;
	#10 counter$count = 88950;
	#10 counter$count = 88951;
	#10 counter$count = 88952;
	#10 counter$count = 88953;
	#10 counter$count = 88954;
	#10 counter$count = 88955;
	#10 counter$count = 88956;
	#10 counter$count = 88957;
	#10 counter$count = 88958;
	#10 counter$count = 88959;
	#10 counter$count = 88960;
	#10 counter$count = 88961;
	#10 counter$count = 88962;
	#10 counter$count = 88963;
	#10 counter$count = 88964;
	#10 counter$count = 88965;
	#10 counter$count = 88966;
	#10 counter$count = 88967;
	#10 counter$count = 88968;
	#10 counter$count = 88969;
	#10 counter$count = 88970;
	#10 counter$count = 88971;
	#10 counter$count = 88972;
	#10 counter$count = 88973;
	#10 counter$count = 88974;
	#10 counter$count = 88975;
	#10 counter$count = 88976;
	#10 counter$count = 88977;
	#10 counter$count = 88978;
	#10 counter$count = 88979;
	#10 counter$count = 88980;
	#10 counter$count = 88981;
	#10 counter$count = 88982;
	#10 counter$count = 88983;
	#10 counter$count = 88984;
	#10 counter$count = 88985;
	#10 counter$count = 88986;
	#10 counter$count = 88987;
	#10 counter$count = 88988;
	#10 counter$count = 88989;
	#10 counter$count = 88990;
	#10 counter$count = 88991;
	#10 counter$count = 88992;
	#10 counter$count = 88993;
	#10 counter$count = 88994;
	#10 counter$count = 88995;
	#10 counter$count = 88996;
	#10 counter$count = 88997;
	#10 counter$count = 88998;
	#10 counter$count = 88999;
	#10 counter$count = 89000;
	#10 counter$count = 89001;
	#10 counter$count = 89002;
	#10 counter$count = 89003;
	#10 counter$count = 89004;
	#10 counter$count = 89005;
	#10 counter$count = 89006;
	#10 counter$count = 89007;
	#10 counter$count = 89008;
	#10 counter$count = 89009;
	#10 counter$count = 89010;
	#10 counter$count = 89011;
	#10 counter$count = 89012;
	#10 counter$count = 89013;
	#10 counter$count = 89014;
	#10 counter$count = 89015;
	#10 counter$count = 89016;
	#10 counter$count = 89017;
	#10 counter$count = 89018;
	#10 counter$count = 89019;
	#10 counter$count = 89020;
	#10 counter$count = 89021;
	#10 counter$count = 89022;
	#10 counter$count = 89023;
	#10 counter$count = 89024;
	#10 counter$count = 89025;
	#10 counter$count = 89026;
	#10 counter$count = 89027;
	#10 counter$count = 89028;
	#10 counter$count = 89029;
	#10 counter$count = 89030;
	#10 counter$count = 89031;
	#10 counter$count = 89032;
	#10 counter$count = 89033;
	#10 counter$count = 89034;
	#10 counter$count = 89035;
	#10 counter$count = 89036;
	#10 counter$count = 89037;
	#10 counter$count = 89038;
	#10 counter$count = 89039;
	#10 counter$count = 89040;
	#10 counter$count = 89041;
	#10 counter$count = 89042;
	#10 counter$count = 89043;
	#10 counter$count = 89044;
	#10 counter$count = 89045;
	#10 counter$count = 89046;
	#10 counter$count = 89047;
	#10 counter$count = 89048;
	#10 counter$count = 89049;
	#10 counter$count = 89050;
	#10 counter$count = 89051;
	#10 counter$count = 89052;
	#10 counter$count = 89053;
	#10 counter$count = 89054;
	#10 counter$count = 89055;
	#10 counter$count = 89056;
	#10 counter$count = 89057;
	#10 counter$count = 89058;
	#10 counter$count = 89059;
	#10 counter$count = 89060;
	#10 counter$count = 89061;
	#10 counter$count = 89062;
	#10 counter$count = 89063;
	#10 counter$count = 89064;
	#10 counter$count = 89065;
	#10 counter$count = 89066;
	#10 counter$count = 89067;
	#10 counter$count = 89068;
	#10 counter$count = 89069;
	#10 counter$count = 89070;
	#10 counter$count = 89071;
	#10 counter$count = 89072;
	#10 counter$count = 89073;
	#10 counter$count = 89074;
	#10 counter$count = 89075;
	#10 counter$count = 89076;
	#10 counter$count = 89077;
	#10 counter$count = 89078;
	#10 counter$count = 89079;
	#10 counter$count = 89080;
	#10 counter$count = 89081;
	#10 counter$count = 89082;
	#10 counter$count = 89083;
	#10 counter$count = 89084;
	#10 counter$count = 89085;
	#10 counter$count = 89086;
	#10 counter$count = 89087;
	#10 counter$count = 89088;
	#10 counter$count = 89089;
	#10 counter$count = 89090;
	#10 counter$count = 89091;
	#10 counter$count = 89092;
	#10 counter$count = 89093;
	#10 counter$count = 89094;
	#10 counter$count = 89095;
	#10 counter$count = 89096;
	#10 counter$count = 89097;
	#10 counter$count = 89098;
	#10 counter$count = 89099;
	#10 counter$count = 89100;
	#10 counter$count = 89101;
	#10 counter$count = 89102;
	#10 counter$count = 89103;
	#10 counter$count = 89104;
	#10 counter$count = 89105;
	#10 counter$count = 89106;
	#10 counter$count = 89107;
	#10 counter$count = 89108;
	#10 counter$count = 89109;
	#10 counter$count = 89110;
	#10 counter$count = 89111;
	#10 counter$count = 89112;
	#10 counter$count = 89113;
	#10 counter$count = 89114;
	#10 counter$count = 89115;
	#10 counter$count = 89116;
	#10 counter$count = 89117;
	#10 counter$count = 89118;
	#10 counter$count = 89119;
	#10 counter$count = 89120;
	#10 counter$count = 89121;
	#10 counter$count = 89122;
	#10 counter$count = 89123;
	#10 counter$count = 89124;
	#10 counter$count = 89125;
	#10 counter$count = 89126;
	#10 counter$count = 89127;
	#10 counter$count = 89128;
	#10 counter$count = 89129;
	#10 counter$count = 89130;
	#10 counter$count = 89131;
	#10 counter$count = 89132;
	#10 counter$count = 89133;
	#10 counter$count = 89134;
	#10 counter$count = 89135;
	#10 counter$count = 89136;
	#10 counter$count = 89137;
	#10 counter$count = 89138;
	#10 counter$count = 89139;
	#10 counter$count = 89140;
	#10 counter$count = 89141;
	#10 counter$count = 89142;
	#10 counter$count = 89143;
	#10 counter$count = 89144;
	#10 counter$count = 89145;
	#10 counter$count = 89146;
	#10 counter$count = 89147;
	#10 counter$count = 89148;
	#10 counter$count = 89149;
	#10 counter$count = 89150;
	#10 counter$count = 89151;
	#10 counter$count = 89152;
	#10 counter$count = 89153;
	#10 counter$count = 89154;
	#10 counter$count = 89155;
	#10 counter$count = 89156;
	#10 counter$count = 89157;
	#10 counter$count = 89158;
	#10 counter$count = 89159;
	#10 counter$count = 89160;
	#10 counter$count = 89161;
	#10 counter$count = 89162;
	#10 counter$count = 89163;
	#10 counter$count = 89164;
	#10 counter$count = 89165;
	#10 counter$count = 89166;
	#10 counter$count = 89167;
	#10 counter$count = 89168;
	#10 counter$count = 89169;
	#10 counter$count = 89170;
	#10 counter$count = 89171;
	#10 counter$count = 89172;
	#10 counter$count = 89173;
	#10 counter$count = 89174;
	#10 counter$count = 89175;
	#10 counter$count = 89176;
	#10 counter$count = 89177;
	#10 counter$count = 89178;
	#10 counter$count = 89179;
	#10 counter$count = 89180;
	#10 counter$count = 89181;
	#10 counter$count = 89182;
	#10 counter$count = 89183;
	#10 counter$count = 89184;
	#10 counter$count = 89185;
	#10 counter$count = 89186;
	#10 counter$count = 89187;
	#10 counter$count = 89188;
	#10 counter$count = 89189;
	#10 counter$count = 89190;
	#10 counter$count = 89191;
	#10 counter$count = 89192;
	#10 counter$count = 89193;
	#10 counter$count = 89194;
	#10 counter$count = 89195;
	#10 counter$count = 89196;
	#10 counter$count = 89197;
	#10 counter$count = 89198;
	#10 counter$count = 89199;
	#10 counter$count = 89200;
	#10 counter$count = 89201;
	#10 counter$count = 89202;
	#10 counter$count = 89203;
	#10 counter$count = 89204;
	#10 counter$count = 89205;
	#10 counter$count = 89206;
	#10 counter$count = 89207;
	#10 counter$count = 89208;
	#10 counter$count = 89209;
	#10 counter$count = 89210;
	#10 counter$count = 89211;
	#10 counter$count = 89212;
	#10 counter$count = 89213;
	#10 counter$count = 89214;
	#10 counter$count = 89215;
	#10 counter$count = 89216;
	#10 counter$count = 89217;
	#10 counter$count = 89218;
	#10 counter$count = 89219;
	#10 counter$count = 89220;
	#10 counter$count = 89221;
	#10 counter$count = 89222;
	#10 counter$count = 89223;
	#10 counter$count = 89224;
	#10 counter$count = 89225;
	#10 counter$count = 89226;
	#10 counter$count = 89227;
	#10 counter$count = 89228;
	#10 counter$count = 89229;
	#10 counter$count = 89230;
	#10 counter$count = 89231;
	#10 counter$count = 89232;
	#10 counter$count = 89233;
	#10 counter$count = 89234;
	#10 counter$count = 89235;
	#10 counter$count = 89236;
	#10 counter$count = 89237;
	#10 counter$count = 89238;
	#10 counter$count = 89239;
	#10 counter$count = 89240;
	#10 counter$count = 89241;
	#10 counter$count = 89242;
	#10 counter$count = 89243;
	#10 counter$count = 89244;
	#10 counter$count = 89245;
	#10 counter$count = 89246;
	#10 counter$count = 89247;
	#10 counter$count = 89248;
	#10 counter$count = 89249;
	#10 counter$count = 89250;
	#10 counter$count = 89251;
	#10 counter$count = 89252;
	#10 counter$count = 89253;
	#10 counter$count = 89254;
	#10 counter$count = 89255;
	#10 counter$count = 89256;
	#10 counter$count = 89257;
	#10 counter$count = 89258;
	#10 counter$count = 89259;
	#10 counter$count = 89260;
	#10 counter$count = 89261;
	#10 counter$count = 89262;
	#10 counter$count = 89263;
	#10 counter$count = 89264;
	#10 counter$count = 89265;
	#10 counter$count = 89266;
	#10 counter$count = 89267;
	#10 counter$count = 89268;
	#10 counter$count = 89269;
	#10 counter$count = 89270;
	#10 counter$count = 89271;
	#10 counter$count = 89272;
	#10 counter$count = 89273;
	#10 counter$count = 89274;
	#10 counter$count = 89275;
	#10 counter$count = 89276;
	#10 counter$count = 89277;
	#10 counter$count = 89278;
	#10 counter$count = 89279;
	#10 counter$count = 89280;
	#10 counter$count = 89281;
	#10 counter$count = 89282;
	#10 counter$count = 89283;
	#10 counter$count = 89284;
	#10 counter$count = 89285;
	#10 counter$count = 89286;
	#10 counter$count = 89287;
	#10 counter$count = 89288;
	#10 counter$count = 89289;
	#10 counter$count = 89290;
	#10 counter$count = 89291;
	#10 counter$count = 89292;
	#10 counter$count = 89293;
	#10 counter$count = 89294;
	#10 counter$count = 89295;
	#10 counter$count = 89296;
	#10 counter$count = 89297;
	#10 counter$count = 89298;
	#10 counter$count = 89299;
	#10 counter$count = 89300;
	#10 counter$count = 89301;
	#10 counter$count = 89302;
	#10 counter$count = 89303;
	#10 counter$count = 89304;
	#10 counter$count = 89305;
	#10 counter$count = 89306;
	#10 counter$count = 89307;
	#10 counter$count = 89308;
	#10 counter$count = 89309;
	#10 counter$count = 89310;
	#10 counter$count = 89311;
	#10 counter$count = 89312;
	#10 counter$count = 89313;
	#10 counter$count = 89314;
	#10 counter$count = 89315;
	#10 counter$count = 89316;
	#10 counter$count = 89317;
	#10 counter$count = 89318;
	#10 counter$count = 89319;
	#10 counter$count = 89320;
	#10 counter$count = 89321;
	#10 counter$count = 89322;
	#10 counter$count = 89323;
	#10 counter$count = 89324;
	#10 counter$count = 89325;
	#10 counter$count = 89326;
	#10 counter$count = 89327;
	#10 counter$count = 89328;
	#10 counter$count = 89329;
	#10 counter$count = 89330;
	#10 counter$count = 89331;
	#10 counter$count = 89332;
	#10 counter$count = 89333;
	#10 counter$count = 89334;
	#10 counter$count = 89335;
	#10 counter$count = 89336;
	#10 counter$count = 89337;
	#10 counter$count = 89338;
	#10 counter$count = 89339;
	#10 counter$count = 89340;
	#10 counter$count = 89341;
	#10 counter$count = 89342;
	#10 counter$count = 89343;
	#10 counter$count = 89344;
	#10 counter$count = 89345;
	#10 counter$count = 89346;
	#10 counter$count = 89347;
	#10 counter$count = 89348;
	#10 counter$count = 89349;
	#10 counter$count = 89350;
	#10 counter$count = 89351;
	#10 counter$count = 89352;
	#10 counter$count = 89353;
	#10 counter$count = 89354;
	#10 counter$count = 89355;
	#10 counter$count = 89356;
	#10 counter$count = 89357;
	#10 counter$count = 89358;
	#10 counter$count = 89359;
	#10 counter$count = 89360;
	#10 counter$count = 89361;
	#10 counter$count = 89362;
	#10 counter$count = 89363;
	#10 counter$count = 89364;
	#10 counter$count = 89365;
	#10 counter$count = 89366;
	#10 counter$count = 89367;
	#10 counter$count = 89368;
	#10 counter$count = 89369;
	#10 counter$count = 89370;
	#10 counter$count = 89371;
	#10 counter$count = 89372;
	#10 counter$count = 89373;
	#10 counter$count = 89374;
	#10 counter$count = 89375;
	#10 counter$count = 89376;
	#10 counter$count = 89377;
	#10 counter$count = 89378;
	#10 counter$count = 89379;
	#10 counter$count = 89380;
	#10 counter$count = 89381;
	#10 counter$count = 89382;
	#10 counter$count = 89383;
	#10 counter$count = 89384;
	#10 counter$count = 89385;
	#10 counter$count = 89386;
	#10 counter$count = 89387;
	#10 counter$count = 89388;
	#10 counter$count = 89389;
	#10 counter$count = 89390;
	#10 counter$count = 89391;
	#10 counter$count = 89392;
	#10 counter$count = 89393;
	#10 counter$count = 89394;
	#10 counter$count = 89395;
	#10 counter$count = 89396;
	#10 counter$count = 89397;
	#10 counter$count = 89398;
	#10 counter$count = 89399;
	#10 counter$count = 89400;
	#10 counter$count = 89401;
	#10 counter$count = 89402;
	#10 counter$count = 89403;
	#10 counter$count = 89404;
	#10 counter$count = 89405;
	#10 counter$count = 89406;
	#10 counter$count = 89407;
	#10 counter$count = 89408;
	#10 counter$count = 89409;
	#10 counter$count = 89410;
	#10 counter$count = 89411;
	#10 counter$count = 89412;
	#10 counter$count = 89413;
	#10 counter$count = 89414;
	#10 counter$count = 89415;
	#10 counter$count = 89416;
	#10 counter$count = 89417;
	#10 counter$count = 89418;
	#10 counter$count = 89419;
	#10 counter$count = 89420;
	#10 counter$count = 89421;
	#10 counter$count = 89422;
	#10 counter$count = 89423;
	#10 counter$count = 89424;
	#10 counter$count = 89425;
	#10 counter$count = 89426;
	#10 counter$count = 89427;
	#10 counter$count = 89428;
	#10 counter$count = 89429;
	#10 counter$count = 89430;
	#10 counter$count = 89431;
	#10 counter$count = 89432;
	#10 counter$count = 89433;
	#10 counter$count = 89434;
	#10 counter$count = 89435;
	#10 counter$count = 89436;
	#10 counter$count = 89437;
	#10 counter$count = 89438;
	#10 counter$count = 89439;
	#10 counter$count = 89440;
	#10 counter$count = 89441;
	#10 counter$count = 89442;
	#10 counter$count = 89443;
	#10 counter$count = 89444;
	#10 counter$count = 89445;
	#10 counter$count = 89446;
	#10 counter$count = 89447;
	#10 counter$count = 89448;
	#10 counter$count = 89449;
	#10 counter$count = 89450;
	#10 counter$count = 89451;
	#10 counter$count = 89452;
	#10 counter$count = 89453;
	#10 counter$count = 89454;
	#10 counter$count = 89455;
	#10 counter$count = 89456;
	#10 counter$count = 89457;
	#10 counter$count = 89458;
	#10 counter$count = 89459;
	#10 counter$count = 89460;
	#10 counter$count = 89461;
	#10 counter$count = 89462;
	#10 counter$count = 89463;
	#10 counter$count = 89464;
	#10 counter$count = 89465;
	#10 counter$count = 89466;
	#10 counter$count = 89467;
	#10 counter$count = 89468;
	#10 counter$count = 89469;
	#10 counter$count = 89470;
	#10 counter$count = 89471;
	#10 counter$count = 89472;
	#10 counter$count = 89473;
	#10 counter$count = 89474;
	#10 counter$count = 89475;
	#10 counter$count = 89476;
	#10 counter$count = 89477;
	#10 counter$count = 89478;
	#10 counter$count = 89479;
	#10 counter$count = 89480;
	#10 counter$count = 89481;
	#10 counter$count = 89482;
	#10 counter$count = 89483;
	#10 counter$count = 89484;
	#10 counter$count = 89485;
	#10 counter$count = 89486;
	#10 counter$count = 89487;
	#10 counter$count = 89488;
	#10 counter$count = 89489;
	#10 counter$count = 89490;
	#10 counter$count = 89491;
	#10 counter$count = 89492;
	#10 counter$count = 89493;
	#10 counter$count = 89494;
	#10 counter$count = 89495;
	#10 counter$count = 89496;
	#10 counter$count = 89497;
	#10 counter$count = 89498;
	#10 counter$count = 89499;
	#10 counter$count = 89500;
	#10 counter$count = 89501;
	#10 counter$count = 89502;
	#10 counter$count = 89503;
	#10 counter$count = 89504;
	#10 counter$count = 89505;
	#10 counter$count = 89506;
	#10 counter$count = 89507;
	#10 counter$count = 89508;
	#10 counter$count = 89509;
	#10 counter$count = 89510;
	#10 counter$count = 89511;
	#10 counter$count = 89512;
	#10 counter$count = 89513;
	#10 counter$count = 89514;
	#10 counter$count = 89515;
	#10 counter$count = 89516;
	#10 counter$count = 89517;
	#10 counter$count = 89518;
	#10 counter$count = 89519;
	#10 counter$count = 89520;
	#10 counter$count = 89521;
	#10 counter$count = 89522;
	#10 counter$count = 89523;
	#10 counter$count = 89524;
	#10 counter$count = 89525;
	#10 counter$count = 89526;
	#10 counter$count = 89527;
	#10 counter$count = 89528;
	#10 counter$count = 89529;
	#10 counter$count = 89530;
	#10 counter$count = 89531;
	#10 counter$count = 89532;
	#10 counter$count = 89533;
	#10 counter$count = 89534;
	#10 counter$count = 89535;
	#10 counter$count = 89536;
	#10 counter$count = 89537;
	#10 counter$count = 89538;
	#10 counter$count = 89539;
	#10 counter$count = 89540;
	#10 counter$count = 89541;
	#10 counter$count = 89542;
	#10 counter$count = 89543;
	#10 counter$count = 89544;
	#10 counter$count = 89545;
	#10 counter$count = 89546;
	#10 counter$count = 89547;
	#10 counter$count = 89548;
	#10 counter$count = 89549;
	#10 counter$count = 89550;
	#10 counter$count = 89551;
	#10 counter$count = 89552;
	#10 counter$count = 89553;
	#10 counter$count = 89554;
	#10 counter$count = 89555;
	#10 counter$count = 89556;
	#10 counter$count = 89557;
	#10 counter$count = 89558;
	#10 counter$count = 89559;
	#10 counter$count = 89560;
	#10 counter$count = 89561;
	#10 counter$count = 89562;
	#10 counter$count = 89563;
	#10 counter$count = 89564;
	#10 counter$count = 89565;
	#10 counter$count = 89566;
	#10 counter$count = 89567;
	#10 counter$count = 89568;
	#10 counter$count = 89569;
	#10 counter$count = 89570;
	#10 counter$count = 89571;
	#10 counter$count = 89572;
	#10 counter$count = 89573;
	#10 counter$count = 89574;
	#10 counter$count = 89575;
	#10 counter$count = 89576;
	#10 counter$count = 89577;
	#10 counter$count = 89578;
	#10 counter$count = 89579;
	#10 counter$count = 89580;
	#10 counter$count = 89581;
	#10 counter$count = 89582;
	#10 counter$count = 89583;
	#10 counter$count = 89584;
	#10 counter$count = 89585;
	#10 counter$count = 89586;
	#10 counter$count = 89587;
	#10 counter$count = 89588;
	#10 counter$count = 89589;
	#10 counter$count = 89590;
	#10 counter$count = 89591;
	#10 counter$count = 89592;
	#10 counter$count = 89593;
	#10 counter$count = 89594;
	#10 counter$count = 89595;
	#10 counter$count = 89596;
	#10 counter$count = 89597;
	#10 counter$count = 89598;
	#10 counter$count = 89599;
	#10 counter$count = 89600;
	#10 counter$count = 89601;
	#10 counter$count = 89602;
	#10 counter$count = 89603;
	#10 counter$count = 89604;
	#10 counter$count = 89605;
	#10 counter$count = 89606;
	#10 counter$count = 89607;
	#10 counter$count = 89608;
	#10 counter$count = 89609;
	#10 counter$count = 89610;
	#10 counter$count = 89611;
	#10 counter$count = 89612;
	#10 counter$count = 89613;
	#10 counter$count = 89614;
	#10 counter$count = 89615;
	#10 counter$count = 89616;
	#10 counter$count = 89617;
	#10 counter$count = 89618;
	#10 counter$count = 89619;
	#10 counter$count = 89620;
	#10 counter$count = 89621;
	#10 counter$count = 89622;
	#10 counter$count = 89623;
	#10 counter$count = 89624;
	#10 counter$count = 89625;
	#10 counter$count = 89626;
	#10 counter$count = 89627;
	#10 counter$count = 89628;
	#10 counter$count = 89629;
	#10 counter$count = 89630;
	#10 counter$count = 89631;
	#10 counter$count = 89632;
	#10 counter$count = 89633;
	#10 counter$count = 89634;
	#10 counter$count = 89635;
	#10 counter$count = 89636;
	#10 counter$count = 89637;
	#10 counter$count = 89638;
	#10 counter$count = 89639;
	#10 counter$count = 89640;
	#10 counter$count = 89641;
	#10 counter$count = 89642;
	#10 counter$count = 89643;
	#10 counter$count = 89644;
	#10 counter$count = 89645;
	#10 counter$count = 89646;
	#10 counter$count = 89647;
	#10 counter$count = 89648;
	#10 counter$count = 89649;
	#10 counter$count = 89650;
	#10 counter$count = 89651;
	#10 counter$count = 89652;
	#10 counter$count = 89653;
	#10 counter$count = 89654;
	#10 counter$count = 89655;
	#10 counter$count = 89656;
	#10 counter$count = 89657;
	#10 counter$count = 89658;
	#10 counter$count = 89659;
	#10 counter$count = 89660;
	#10 counter$count = 89661;
	#10 counter$count = 89662;
	#10 counter$count = 89663;
	#10 counter$count = 89664;
	#10 counter$count = 89665;
	#10 counter$count = 89666;
	#10 counter$count = 89667;
	#10 counter$count = 89668;
	#10 counter$count = 89669;
	#10 counter$count = 89670;
	#10 counter$count = 89671;
	#10 counter$count = 89672;
	#10 counter$count = 89673;
	#10 counter$count = 89674;
	#10 counter$count = 89675;
	#10 counter$count = 89676;
	#10 counter$count = 89677;
	#10 counter$count = 89678;
	#10 counter$count = 89679;
	#10 counter$count = 89680;
	#10 counter$count = 89681;
	#10 counter$count = 89682;
	#10 counter$count = 89683;
	#10 counter$count = 89684;
	#10 counter$count = 89685;
	#10 counter$count = 89686;
	#10 counter$count = 89687;
	#10 counter$count = 89688;
	#10 counter$count = 89689;
	#10 counter$count = 89690;
	#10 counter$count = 89691;
	#10 counter$count = 89692;
	#10 counter$count = 89693;
	#10 counter$count = 89694;
	#10 counter$count = 89695;
	#10 counter$count = 89696;
	#10 counter$count = 89697;
	#10 counter$count = 89698;
	#10 counter$count = 89699;
	#10 counter$count = 89700;
	#10 counter$count = 89701;
	#10 counter$count = 89702;
	#10 counter$count = 89703;
	#10 counter$count = 89704;
	#10 counter$count = 89705;
	#10 counter$count = 89706;
	#10 counter$count = 89707;
	#10 counter$count = 89708;
	#10 counter$count = 89709;
	#10 counter$count = 89710;
	#10 counter$count = 89711;
	#10 counter$count = 89712;
	#10 counter$count = 89713;
	#10 counter$count = 89714;
	#10 counter$count = 89715;
	#10 counter$count = 89716;
	#10 counter$count = 89717;
	#10 counter$count = 89718;
	#10 counter$count = 89719;
	#10 counter$count = 89720;
	#10 counter$count = 89721;
	#10 counter$count = 89722;
	#10 counter$count = 89723;
	#10 counter$count = 89724;
	#10 counter$count = 89725;
	#10 counter$count = 89726;
	#10 counter$count = 89727;
	#10 counter$count = 89728;
	#10 counter$count = 89729;
	#10 counter$count = 89730;
	#10 counter$count = 89731;
	#10 counter$count = 89732;
	#10 counter$count = 89733;
	#10 counter$count = 89734;
	#10 counter$count = 89735;
	#10 counter$count = 89736;
	#10 counter$count = 89737;
	#10 counter$count = 89738;
	#10 counter$count = 89739;
	#10 counter$count = 89740;
	#10 counter$count = 89741;
	#10 counter$count = 89742;
	#10 counter$count = 89743;
	#10 counter$count = 89744;
	#10 counter$count = 89745;
	#10 counter$count = 89746;
	#10 counter$count = 89747;
	#10 counter$count = 89748;
	#10 counter$count = 89749;
	#10 counter$count = 89750;
	#10 counter$count = 89751;
	#10 counter$count = 89752;
	#10 counter$count = 89753;
	#10 counter$count = 89754;
	#10 counter$count = 89755;
	#10 counter$count = 89756;
	#10 counter$count = 89757;
	#10 counter$count = 89758;
	#10 counter$count = 89759;
	#10 counter$count = 89760;
	#10 counter$count = 89761;
	#10 counter$count = 89762;
	#10 counter$count = 89763;
	#10 counter$count = 89764;
	#10 counter$count = 89765;
	#10 counter$count = 89766;
	#10 counter$count = 89767;
	#10 counter$count = 89768;
	#10 counter$count = 89769;
	#10 counter$count = 89770;
	#10 counter$count = 89771;
	#10 counter$count = 89772;
	#10 counter$count = 89773;
	#10 counter$count = 89774;
	#10 counter$count = 89775;
	#10 counter$count = 89776;
	#10 counter$count = 89777;
	#10 counter$count = 89778;
	#10 counter$count = 89779;
	#10 counter$count = 89780;
	#10 counter$count = 89781;
	#10 counter$count = 89782;
	#10 counter$count = 89783;
	#10 counter$count = 89784;
	#10 counter$count = 89785;
	#10 counter$count = 89786;
	#10 counter$count = 89787;
	#10 counter$count = 89788;
	#10 counter$count = 89789;
	#10 counter$count = 89790;
	#10 counter$count = 89791;
	#10 counter$count = 89792;
	#10 counter$count = 89793;
	#10 counter$count = 89794;
	#10 counter$count = 89795;
	#10 counter$count = 89796;
	#10 counter$count = 89797;
	#10 counter$count = 89798;
	#10 counter$count = 89799;
	#10 counter$count = 89800;
	#10 counter$count = 89801;
	#10 counter$count = 89802;
	#10 counter$count = 89803;
	#10 counter$count = 89804;
	#10 counter$count = 89805;
	#10 counter$count = 89806;
	#10 counter$count = 89807;
	#10 counter$count = 89808;
	#10 counter$count = 89809;
	#10 counter$count = 89810;
	#10 counter$count = 89811;
	#10 counter$count = 89812;
	#10 counter$count = 89813;
	#10 counter$count = 89814;
	#10 counter$count = 89815;
	#10 counter$count = 89816;
	#10 counter$count = 89817;
	#10 counter$count = 89818;
	#10 counter$count = 89819;
	#10 counter$count = 89820;
	#10 counter$count = 89821;
	#10 counter$count = 89822;
	#10 counter$count = 89823;
	#10 counter$count = 89824;
	#10 counter$count = 89825;
	#10 counter$count = 89826;
	#10 counter$count = 89827;
	#10 counter$count = 89828;
	#10 counter$count = 89829;
	#10 counter$count = 89830;
	#10 counter$count = 89831;
	#10 counter$count = 89832;
	#10 counter$count = 89833;
	#10 counter$count = 89834;
	#10 counter$count = 89835;
	#10 counter$count = 89836;
	#10 counter$count = 89837;
	#10 counter$count = 89838;
	#10 counter$count = 89839;
	#10 counter$count = 89840;
	#10 counter$count = 89841;
	#10 counter$count = 89842;
	#10 counter$count = 89843;
	#10 counter$count = 89844;
	#10 counter$count = 89845;
	#10 counter$count = 89846;
	#10 counter$count = 89847;
	#10 counter$count = 89848;
	#10 counter$count = 89849;
	#10 counter$count = 89850;
	#10 counter$count = 89851;
	#10 counter$count = 89852;
	#10 counter$count = 89853;
	#10 counter$count = 89854;
	#10 counter$count = 89855;
	#10 counter$count = 89856;
	#10 counter$count = 89857;
	#10 counter$count = 89858;
	#10 counter$count = 89859;
	#10 counter$count = 89860;
	#10 counter$count = 89861;
	#10 counter$count = 89862;
	#10 counter$count = 89863;
	#10 counter$count = 89864;
	#10 counter$count = 89865;
	#10 counter$count = 89866;
	#10 counter$count = 89867;
	#10 counter$count = 89868;
	#10 counter$count = 89869;
	#10 counter$count = 89870;
	#10 counter$count = 89871;
	#10 counter$count = 89872;
	#10 counter$count = 89873;
	#10 counter$count = 89874;
	#10 counter$count = 89875;
	#10 counter$count = 89876;
	#10 counter$count = 89877;
	#10 counter$count = 89878;
	#10 counter$count = 89879;
	#10 counter$count = 89880;
	#10 counter$count = 89881;
	#10 counter$count = 89882;
	#10 counter$count = 89883;
	#10 counter$count = 89884;
	#10 counter$count = 89885;
	#10 counter$count = 89886;
	#10 counter$count = 89887;
	#10 counter$count = 89888;
	#10 counter$count = 89889;
	#10 counter$count = 89890;
	#10 counter$count = 89891;
	#10 counter$count = 89892;
	#10 counter$count = 89893;
	#10 counter$count = 89894;
	#10 counter$count = 89895;
	#10 counter$count = 89896;
	#10 counter$count = 89897;
	#10 counter$count = 89898;
	#10 counter$count = 89899;
	#10 counter$count = 89900;
	#10 counter$count = 89901;
	#10 counter$count = 89902;
	#10 counter$count = 89903;
	#10 counter$count = 89904;
	#10 counter$count = 89905;
	#10 counter$count = 89906;
	#10 counter$count = 89907;
	#10 counter$count = 89908;
	#10 counter$count = 89909;
	#10 counter$count = 89910;
	#10 counter$count = 89911;
	#10 counter$count = 89912;
	#10 counter$count = 89913;
	#10 counter$count = 89914;
	#10 counter$count = 89915;
	#10 counter$count = 89916;
	#10 counter$count = 89917;
	#10 counter$count = 89918;
	#10 counter$count = 89919;
	#10 counter$count = 89920;
	#10 counter$count = 89921;
	#10 counter$count = 89922;
	#10 counter$count = 89923;
	#10 counter$count = 89924;
	#10 counter$count = 89925;
	#10 counter$count = 89926;
	#10 counter$count = 89927;
	#10 counter$count = 89928;
	#10 counter$count = 89929;
	#10 counter$count = 89930;
	#10 counter$count = 89931;
	#10 counter$count = 89932;
	#10 counter$count = 89933;
	#10 counter$count = 89934;
	#10 counter$count = 89935;
	#10 counter$count = 89936;
	#10 counter$count = 89937;
	#10 counter$count = 89938;
	#10 counter$count = 89939;
	#10 counter$count = 89940;
	#10 counter$count = 89941;
	#10 counter$count = 89942;
	#10 counter$count = 89943;
	#10 counter$count = 89944;
	#10 counter$count = 89945;
	#10 counter$count = 89946;
	#10 counter$count = 89947;
	#10 counter$count = 89948;
	#10 counter$count = 89949;
	#10 counter$count = 89950;
	#10 counter$count = 89951;
	#10 counter$count = 89952;
	#10 counter$count = 89953;
	#10 counter$count = 89954;
	#10 counter$count = 89955;
	#10 counter$count = 89956;
	#10 counter$count = 89957;
	#10 counter$count = 89958;
	#10 counter$count = 89959;
	#10 counter$count = 89960;
	#10 counter$count = 89961;
	#10 counter$count = 89962;
	#10 counter$count = 89963;
	#10 counter$count = 89964;
	#10 counter$count = 89965;
	#10 counter$count = 89966;
	#10 counter$count = 89967;
	#10 counter$count = 89968;
	#10 counter$count = 89969;
	#10 counter$count = 89970;
	#10 counter$count = 89971;
	#10 counter$count = 89972;
	#10 counter$count = 89973;
	#10 counter$count = 89974;
	#10 counter$count = 89975;
	#10 counter$count = 89976;
	#10 counter$count = 89977;
	#10 counter$count = 89978;
	#10 counter$count = 89979;
	#10 counter$count = 89980;
	#10 counter$count = 89981;
	#10 counter$count = 89982;
	#10 counter$count = 89983;
	#10 counter$count = 89984;
	#10 counter$count = 89985;
	#10 counter$count = 89986;
	#10 counter$count = 89987;
	#10 counter$count = 89988;
	#10 counter$count = 89989;
	#10 counter$count = 89990;
	#10 counter$count = 89991;
	#10 counter$count = 89992;
	#10 counter$count = 89993;
	#10 counter$count = 89994;
	#10 counter$count = 89995;
	#10 counter$count = 89996;
	#10 counter$count = 89997;
	#10 counter$count = 89998;
	#10 counter$count = 89999;
	#10 counter$count = 90000;
	#10 counter$count = 90001;
	#10 counter$count = 90002;
	#10 counter$count = 90003;
	#10 counter$count = 90004;
	#10 counter$count = 90005;
	#10 counter$count = 90006;
	#10 counter$count = 90007;
	#10 counter$count = 90008;
	#10 counter$count = 90009;
	#10 counter$count = 90010;
	#10 counter$count = 90011;
	#10 counter$count = 90012;
	#10 counter$count = 90013;
	#10 counter$count = 90014;
	#10 counter$count = 90015;
	#10 counter$count = 90016;
	#10 counter$count = 90017;
	#10 counter$count = 90018;
	#10 counter$count = 90019;
	#10 counter$count = 90020;
	#10 counter$count = 90021;
	#10 counter$count = 90022;
	#10 counter$count = 90023;
	#10 counter$count = 90024;
	#10 counter$count = 90025;
	#10 counter$count = 90026;
	#10 counter$count = 90027;
	#10 counter$count = 90028;
	#10 counter$count = 90029;
	#10 counter$count = 90030;
	#10 counter$count = 90031;
	#10 counter$count = 90032;
	#10 counter$count = 90033;
	#10 counter$count = 90034;
	#10 counter$count = 90035;
	#10 counter$count = 90036;
	#10 counter$count = 90037;
	#10 counter$count = 90038;
	#10 counter$count = 90039;
	#10 counter$count = 90040;
	#10 counter$count = 90041;
	#10 counter$count = 90042;
	#10 counter$count = 90043;
	#10 counter$count = 90044;
	#10 counter$count = 90045;
	#10 counter$count = 90046;
	#10 counter$count = 90047;
	#10 counter$count = 90048;
	#10 counter$count = 90049;
	#10 counter$count = 90050;
	#10 counter$count = 90051;
	#10 counter$count = 90052;
	#10 counter$count = 90053;
	#10 counter$count = 90054;
	#10 counter$count = 90055;
	#10 counter$count = 90056;
	#10 counter$count = 90057;
	#10 counter$count = 90058;
	#10 counter$count = 90059;
	#10 counter$count = 90060;
	#10 counter$count = 90061;
	#10 counter$count = 90062;
	#10 counter$count = 90063;
	#10 counter$count = 90064;
	#10 counter$count = 90065;
	#10 counter$count = 90066;
	#10 counter$count = 90067;
	#10 counter$count = 90068;
	#10 counter$count = 90069;
	#10 counter$count = 90070;
	#10 counter$count = 90071;
	#10 counter$count = 90072;
	#10 counter$count = 90073;
	#10 counter$count = 90074;
	#10 counter$count = 90075;
	#10 counter$count = 90076;
	#10 counter$count = 90077;
	#10 counter$count = 90078;
	#10 counter$count = 90079;
	#10 counter$count = 90080;
	#10 counter$count = 90081;
	#10 counter$count = 90082;
	#10 counter$count = 90083;
	#10 counter$count = 90084;
	#10 counter$count = 90085;
	#10 counter$count = 90086;
	#10 counter$count = 90087;
	#10 counter$count = 90088;
	#10 counter$count = 90089;
	#10 counter$count = 90090;
	#10 counter$count = 90091;
	#10 counter$count = 90092;
	#10 counter$count = 90093;
	#10 counter$count = 90094;
	#10 counter$count = 90095;
	#10 counter$count = 90096;
	#10 counter$count = 90097;
	#10 counter$count = 90098;
	#10 counter$count = 90099;
	#10 counter$count = 90100;
	#10 counter$count = 90101;
	#10 counter$count = 90102;
	#10 counter$count = 90103;
	#10 counter$count = 90104;
	#10 counter$count = 90105;
	#10 counter$count = 90106;
	#10 counter$count = 90107;
	#10 counter$count = 90108;
	#10 counter$count = 90109;
	#10 counter$count = 90110;
	#10 counter$count = 90111;
	#10 counter$count = 90112;
	#10 counter$count = 90113;
	#10 counter$count = 90114;
	#10 counter$count = 90115;
	#10 counter$count = 90116;
	#10 counter$count = 90117;
	#10 counter$count = 90118;
	#10 counter$count = 90119;
	#10 counter$count = 90120;
	#10 counter$count = 90121;
	#10 counter$count = 90122;
	#10 counter$count = 90123;
	#10 counter$count = 90124;
	#10 counter$count = 90125;
	#10 counter$count = 90126;
	#10 counter$count = 90127;
	#10 counter$count = 90128;
	#10 counter$count = 90129;
	#10 counter$count = 90130;
	#10 counter$count = 90131;
	#10 counter$count = 90132;
	#10 counter$count = 90133;
	#10 counter$count = 90134;
	#10 counter$count = 90135;
	#10 counter$count = 90136;
	#10 counter$count = 90137;
	#10 counter$count = 90138;
	#10 counter$count = 90139;
	#10 counter$count = 90140;
	#10 counter$count = 90141;
	#10 counter$count = 90142;
	#10 counter$count = 90143;
	#10 counter$count = 90144;
	#10 counter$count = 90145;
	#10 counter$count = 90146;
	#10 counter$count = 90147;
	#10 counter$count = 90148;
	#10 counter$count = 90149;
	#10 counter$count = 90150;
	#10 counter$count = 90151;
	#10 counter$count = 90152;
	#10 counter$count = 90153;
	#10 counter$count = 90154;
	#10 counter$count = 90155;
	#10 counter$count = 90156;
	#10 counter$count = 90157;
	#10 counter$count = 90158;
	#10 counter$count = 90159;
	#10 counter$count = 90160;
	#10 counter$count = 90161;
	#10 counter$count = 90162;
	#10 counter$count = 90163;
	#10 counter$count = 90164;
	#10 counter$count = 90165;
	#10 counter$count = 90166;
	#10 counter$count = 90167;
	#10 counter$count = 90168;
	#10 counter$count = 90169;
	#10 counter$count = 90170;
	#10 counter$count = 90171;
	#10 counter$count = 90172;
	#10 counter$count = 90173;
	#10 counter$count = 90174;
	#10 counter$count = 90175;
	#10 counter$count = 90176;
	#10 counter$count = 90177;
	#10 counter$count = 90178;
	#10 counter$count = 90179;
	#10 counter$count = 90180;
	#10 counter$count = 90181;
	#10 counter$count = 90182;
	#10 counter$count = 90183;
	#10 counter$count = 90184;
	#10 counter$count = 90185;
	#10 counter$count = 90186;
	#10 counter$count = 90187;
	#10 counter$count = 90188;
	#10 counter$count = 90189;
	#10 counter$count = 90190;
	#10 counter$count = 90191;
	#10 counter$count = 90192;
	#10 counter$count = 90193;
	#10 counter$count = 90194;
	#10 counter$count = 90195;
	#10 counter$count = 90196;
	#10 counter$count = 90197;
	#10 counter$count = 90198;
	#10 counter$count = 90199;
	#10 counter$count = 90200;
	#10 counter$count = 90201;
	#10 counter$count = 90202;
	#10 counter$count = 90203;
	#10 counter$count = 90204;
	#10 counter$count = 90205;
	#10 counter$count = 90206;
	#10 counter$count = 90207;
	#10 counter$count = 90208;
	#10 counter$count = 90209;
	#10 counter$count = 90210;
	#10 counter$count = 90211;
	#10 counter$count = 90212;
	#10 counter$count = 90213;
	#10 counter$count = 90214;
	#10 counter$count = 90215;
	#10 counter$count = 90216;
	#10 counter$count = 90217;
	#10 counter$count = 90218;
	#10 counter$count = 90219;
	#10 counter$count = 90220;
	#10 counter$count = 90221;
	#10 counter$count = 90222;
	#10 counter$count = 90223;
	#10 counter$count = 90224;
	#10 counter$count = 90225;
	#10 counter$count = 90226;
	#10 counter$count = 90227;
	#10 counter$count = 90228;
	#10 counter$count = 90229;
	#10 counter$count = 90230;
	#10 counter$count = 90231;
	#10 counter$count = 90232;
	#10 counter$count = 90233;
	#10 counter$count = 90234;
	#10 counter$count = 90235;
	#10 counter$count = 90236;
	#10 counter$count = 90237;
	#10 counter$count = 90238;
	#10 counter$count = 90239;
	#10 counter$count = 90240;
	#10 counter$count = 90241;
	#10 counter$count = 90242;
	#10 counter$count = 90243;
	#10 counter$count = 90244;
	#10 counter$count = 90245;
	#10 counter$count = 90246;
	#10 counter$count = 90247;
	#10 counter$count = 90248;
	#10 counter$count = 90249;
	#10 counter$count = 90250;
	#10 counter$count = 90251;
	#10 counter$count = 90252;
	#10 counter$count = 90253;
	#10 counter$count = 90254;
	#10 counter$count = 90255;
	#10 counter$count = 90256;
	#10 counter$count = 90257;
	#10 counter$count = 90258;
	#10 counter$count = 90259;
	#10 counter$count = 90260;
	#10 counter$count = 90261;
	#10 counter$count = 90262;
	#10 counter$count = 90263;
	#10 counter$count = 90264;
	#10 counter$count = 90265;
	#10 counter$count = 90266;
	#10 counter$count = 90267;
	#10 counter$count = 90268;
	#10 counter$count = 90269;
	#10 counter$count = 90270;
	#10 counter$count = 90271;
	#10 counter$count = 90272;
	#10 counter$count = 90273;
	#10 counter$count = 90274;
	#10 counter$count = 90275;
	#10 counter$count = 90276;
	#10 counter$count = 90277;
	#10 counter$count = 90278;
	#10 counter$count = 90279;
	#10 counter$count = 90280;
	#10 counter$count = 90281;
	#10 counter$count = 90282;
	#10 counter$count = 90283;
	#10 counter$count = 90284;
	#10 counter$count = 90285;
	#10 counter$count = 90286;
	#10 counter$count = 90287;
	#10 counter$count = 90288;
	#10 counter$count = 90289;
	#10 counter$count = 90290;
	#10 counter$count = 90291;
	#10 counter$count = 90292;
	#10 counter$count = 90293;
	#10 counter$count = 90294;
	#10 counter$count = 90295;
	#10 counter$count = 90296;
	#10 counter$count = 90297;
	#10 counter$count = 90298;
	#10 counter$count = 90299;
	#10 counter$count = 90300;
	#10 counter$count = 90301;
	#10 counter$count = 90302;
	#10 counter$count = 90303;
	#10 counter$count = 90304;
	#10 counter$count = 90305;
	#10 counter$count = 90306;
	#10 counter$count = 90307;
	#10 counter$count = 90308;
	#10 counter$count = 90309;
	#10 counter$count = 90310;
	#10 counter$count = 90311;
	#10 counter$count = 90312;
	#10 counter$count = 90313;
	#10 counter$count = 90314;
	#10 counter$count = 90315;
	#10 counter$count = 90316;
	#10 counter$count = 90317;
	#10 counter$count = 90318;
	#10 counter$count = 90319;
	#10 counter$count = 90320;
	#10 counter$count = 90321;
	#10 counter$count = 90322;
	#10 counter$count = 90323;
	#10 counter$count = 90324;
	#10 counter$count = 90325;
	#10 counter$count = 90326;
	#10 counter$count = 90327;
	#10 counter$count = 90328;
	#10 counter$count = 90329;
	#10 counter$count = 90330;
	#10 counter$count = 90331;
	#10 counter$count = 90332;
	#10 counter$count = 90333;
	#10 counter$count = 90334;
	#10 counter$count = 90335;
	#10 counter$count = 90336;
	#10 counter$count = 90337;
	#10 counter$count = 90338;
	#10 counter$count = 90339;
	#10 counter$count = 90340;
	#10 counter$count = 90341;
	#10 counter$count = 90342;
	#10 counter$count = 90343;
	#10 counter$count = 90344;
	#10 counter$count = 90345;
	#10 counter$count = 90346;
	#10 counter$count = 90347;
	#10 counter$count = 90348;
	#10 counter$count = 90349;
	#10 counter$count = 90350;
	#10 counter$count = 90351;
	#10 counter$count = 90352;
	#10 counter$count = 90353;
	#10 counter$count = 90354;
	#10 counter$count = 90355;
	#10 counter$count = 90356;
	#10 counter$count = 90357;
	#10 counter$count = 90358;
	#10 counter$count = 90359;
	#10 counter$count = 90360;
	#10 counter$count = 90361;
	#10 counter$count = 90362;
	#10 counter$count = 90363;
	#10 counter$count = 90364;
	#10 counter$count = 90365;
	#10 counter$count = 90366;
	#10 counter$count = 90367;
	#10 counter$count = 90368;
	#10 counter$count = 90369;
	#10 counter$count = 90370;
	#10 counter$count = 90371;
	#10 counter$count = 90372;
	#10 counter$count = 90373;
	#10 counter$count = 90374;
	#10 counter$count = 90375;
	#10 counter$count = 90376;
	#10 counter$count = 90377;
	#10 counter$count = 90378;
	#10 counter$count = 90379;
	#10 counter$count = 90380;
	#10 counter$count = 90381;
	#10 counter$count = 90382;
	#10 counter$count = 90383;
	#10 counter$count = 90384;
	#10 counter$count = 90385;
	#10 counter$count = 90386;
	#10 counter$count = 90387;
	#10 counter$count = 90388;
	#10 counter$count = 90389;
	#10 counter$count = 90390;
	#10 counter$count = 90391;
	#10 counter$count = 90392;
	#10 counter$count = 90393;
	#10 counter$count = 90394;
	#10 counter$count = 90395;
	#10 counter$count = 90396;
	#10 counter$count = 90397;
	#10 counter$count = 90398;
	#10 counter$count = 90399;
	#10 counter$count = 90400;
	#10 counter$count = 90401;
	#10 counter$count = 90402;
	#10 counter$count = 90403;
	#10 counter$count = 90404;
	#10 counter$count = 90405;
	#10 counter$count = 90406;
	#10 counter$count = 90407;
	#10 counter$count = 90408;
	#10 counter$count = 90409;
	#10 counter$count = 90410;
	#10 counter$count = 90411;
	#10 counter$count = 90412;
	#10 counter$count = 90413;
	#10 counter$count = 90414;
	#10 counter$count = 90415;
	#10 counter$count = 90416;
	#10 counter$count = 90417;
	#10 counter$count = 90418;
	#10 counter$count = 90419;
	#10 counter$count = 90420;
	#10 counter$count = 90421;
	#10 counter$count = 90422;
	#10 counter$count = 90423;
	#10 counter$count = 90424;
	#10 counter$count = 90425;
	#10 counter$count = 90426;
	#10 counter$count = 90427;
	#10 counter$count = 90428;
	#10 counter$count = 90429;
	#10 counter$count = 90430;
	#10 counter$count = 90431;
	#10 counter$count = 90432;
	#10 counter$count = 90433;
	#10 counter$count = 90434;
	#10 counter$count = 90435;
	#10 counter$count = 90436;
	#10 counter$count = 90437;
	#10 counter$count = 90438;
	#10 counter$count = 90439;
	#10 counter$count = 90440;
	#10 counter$count = 90441;
	#10 counter$count = 90442;
	#10 counter$count = 90443;
	#10 counter$count = 90444;
	#10 counter$count = 90445;
	#10 counter$count = 90446;
	#10 counter$count = 90447;
	#10 counter$count = 90448;
	#10 counter$count = 90449;
	#10 counter$count = 90450;
	#10 counter$count = 90451;
	#10 counter$count = 90452;
	#10 counter$count = 90453;
	#10 counter$count = 90454;
	#10 counter$count = 90455;
	#10 counter$count = 90456;
	#10 counter$count = 90457;
	#10 counter$count = 90458;
	#10 counter$count = 90459;
	#10 counter$count = 90460;
	#10 counter$count = 90461;
	#10 counter$count = 90462;
	#10 counter$count = 90463;
	#10 counter$count = 90464;
	#10 counter$count = 90465;
	#10 counter$count = 90466;
	#10 counter$count = 90467;
	#10 counter$count = 90468;
	#10 counter$count = 90469;
	#10 counter$count = 90470;
	#10 counter$count = 90471;
	#10 counter$count = 90472;
	#10 counter$count = 90473;
	#10 counter$count = 90474;
	#10 counter$count = 90475;
	#10 counter$count = 90476;
	#10 counter$count = 90477;
	#10 counter$count = 90478;
	#10 counter$count = 90479;
	#10 counter$count = 90480;
	#10 counter$count = 90481;
	#10 counter$count = 90482;
	#10 counter$count = 90483;
	#10 counter$count = 90484;
	#10 counter$count = 90485;
	#10 counter$count = 90486;
	#10 counter$count = 90487;
	#10 counter$count = 90488;
	#10 counter$count = 90489;
	#10 counter$count = 90490;
	#10 counter$count = 90491;
	#10 counter$count = 90492;
	#10 counter$count = 90493;
	#10 counter$count = 90494;
	#10 counter$count = 90495;
	#10 counter$count = 90496;
	#10 counter$count = 90497;
	#10 counter$count = 90498;
	#10 counter$count = 90499;
	#10 counter$count = 90500;
	#10 counter$count = 90501;
	#10 counter$count = 90502;
	#10 counter$count = 90503;
	#10 counter$count = 90504;
	#10 counter$count = 90505;
	#10 counter$count = 90506;
	#10 counter$count = 90507;
	#10 counter$count = 90508;
	#10 counter$count = 90509;
	#10 counter$count = 90510;
	#10 counter$count = 90511;
	#10 counter$count = 90512;
	#10 counter$count = 90513;
	#10 counter$count = 90514;
	#10 counter$count = 90515;
	#10 counter$count = 90516;
	#10 counter$count = 90517;
	#10 counter$count = 90518;
	#10 counter$count = 90519;
	#10 counter$count = 90520;
	#10 counter$count = 90521;
	#10 counter$count = 90522;
	#10 counter$count = 90523;
	#10 counter$count = 90524;
	#10 counter$count = 90525;
	#10 counter$count = 90526;
	#10 counter$count = 90527;
	#10 counter$count = 90528;
	#10 counter$count = 90529;
	#10 counter$count = 90530;
	#10 counter$count = 90531;
	#10 counter$count = 90532;
	#10 counter$count = 90533;
	#10 counter$count = 90534;
	#10 counter$count = 90535;
	#10 counter$count = 90536;
	#10 counter$count = 90537;
	#10 counter$count = 90538;
	#10 counter$count = 90539;
	#10 counter$count = 90540;
	#10 counter$count = 90541;
	#10 counter$count = 90542;
	#10 counter$count = 90543;
	#10 counter$count = 90544;
	#10 counter$count = 90545;
	#10 counter$count = 90546;
	#10 counter$count = 90547;
	#10 counter$count = 90548;
	#10 counter$count = 90549;
	#10 counter$count = 90550;
	#10 counter$count = 90551;
	#10 counter$count = 90552;
	#10 counter$count = 90553;
	#10 counter$count = 90554;
	#10 counter$count = 90555;
	#10 counter$count = 90556;
	#10 counter$count = 90557;
	#10 counter$count = 90558;
	#10 counter$count = 90559;
	#10 counter$count = 90560;
	#10 counter$count = 90561;
	#10 counter$count = 90562;
	#10 counter$count = 90563;
	#10 counter$count = 90564;
	#10 counter$count = 90565;
	#10 counter$count = 90566;
	#10 counter$count = 90567;
	#10 counter$count = 90568;
	#10 counter$count = 90569;
	#10 counter$count = 90570;
	#10 counter$count = 90571;
	#10 counter$count = 90572;
	#10 counter$count = 90573;
	#10 counter$count = 90574;
	#10 counter$count = 90575;
	#10 counter$count = 90576;
	#10 counter$count = 90577;
	#10 counter$count = 90578;
	#10 counter$count = 90579;
	#10 counter$count = 90580;
	#10 counter$count = 90581;
	#10 counter$count = 90582;
	#10 counter$count = 90583;
	#10 counter$count = 90584;
	#10 counter$count = 90585;
	#10 counter$count = 90586;
	#10 counter$count = 90587;
	#10 counter$count = 90588;
	#10 counter$count = 90589;
	#10 counter$count = 90590;
	#10 counter$count = 90591;
	#10 counter$count = 90592;
	#10 counter$count = 90593;
	#10 counter$count = 90594;
	#10 counter$count = 90595;
	#10 counter$count = 90596;
	#10 counter$count = 90597;
	#10 counter$count = 90598;
	#10 counter$count = 90599;
	#10 counter$count = 90600;
	#10 counter$count = 90601;
	#10 counter$count = 90602;
	#10 counter$count = 90603;
	#10 counter$count = 90604;
	#10 counter$count = 90605;
	#10 counter$count = 90606;
	#10 counter$count = 90607;
	#10 counter$count = 90608;
	#10 counter$count = 90609;
	#10 counter$count = 90610;
	#10 counter$count = 90611;
	#10 counter$count = 90612;
	#10 counter$count = 90613;
	#10 counter$count = 90614;
	#10 counter$count = 90615;
	#10 counter$count = 90616;
	#10 counter$count = 90617;
	#10 counter$count = 90618;
	#10 counter$count = 90619;
	#10 counter$count = 90620;
	#10 counter$count = 90621;
	#10 counter$count = 90622;
	#10 counter$count = 90623;
	#10 counter$count = 90624;
	#10 counter$count = 90625;
	#10 counter$count = 90626;
	#10 counter$count = 90627;
	#10 counter$count = 90628;
	#10 counter$count = 90629;
	#10 counter$count = 90630;
	#10 counter$count = 90631;
	#10 counter$count = 90632;
	#10 counter$count = 90633;
	#10 counter$count = 90634;
	#10 counter$count = 90635;
	#10 counter$count = 90636;
	#10 counter$count = 90637;
	#10 counter$count = 90638;
	#10 counter$count = 90639;
	#10 counter$count = 90640;
	#10 counter$count = 90641;
	#10 counter$count = 90642;
	#10 counter$count = 90643;
	#10 counter$count = 90644;
	#10 counter$count = 90645;
	#10 counter$count = 90646;
	#10 counter$count = 90647;
	#10 counter$count = 90648;
	#10 counter$count = 90649;
	#10 counter$count = 90650;
	#10 counter$count = 90651;
	#10 counter$count = 90652;
	#10 counter$count = 90653;
	#10 counter$count = 90654;
	#10 counter$count = 90655;
	#10 counter$count = 90656;
	#10 counter$count = 90657;
	#10 counter$count = 90658;
	#10 counter$count = 90659;
	#10 counter$count = 90660;
	#10 counter$count = 90661;
	#10 counter$count = 90662;
	#10 counter$count = 90663;
	#10 counter$count = 90664;
	#10 counter$count = 90665;
	#10 counter$count = 90666;
	#10 counter$count = 90667;
	#10 counter$count = 90668;
	#10 counter$count = 90669;
	#10 counter$count = 90670;
	#10 counter$count = 90671;
	#10 counter$count = 90672;
	#10 counter$count = 90673;
	#10 counter$count = 90674;
	#10 counter$count = 90675;
	#10 counter$count = 90676;
	#10 counter$count = 90677;
	#10 counter$count = 90678;
	#10 counter$count = 90679;
	#10 counter$count = 90680;
	#10 counter$count = 90681;
	#10 counter$count = 90682;
	#10 counter$count = 90683;
	#10 counter$count = 90684;
	#10 counter$count = 90685;
	#10 counter$count = 90686;
	#10 counter$count = 90687;
	#10 counter$count = 90688;
	#10 counter$count = 90689;
	#10 counter$count = 90690;
	#10 counter$count = 90691;
	#10 counter$count = 90692;
	#10 counter$count = 90693;
	#10 counter$count = 90694;
	#10 counter$count = 90695;
	#10 counter$count = 90696;
	#10 counter$count = 90697;
	#10 counter$count = 90698;
	#10 counter$count = 90699;
	#10 counter$count = 90700;
	#10 counter$count = 90701;
	#10 counter$count = 90702;
	#10 counter$count = 90703;
	#10 counter$count = 90704;
	#10 counter$count = 90705;
	#10 counter$count = 90706;
	#10 counter$count = 90707;
	#10 counter$count = 90708;
	#10 counter$count = 90709;
	#10 counter$count = 90710;
	#10 counter$count = 90711;
	#10 counter$count = 90712;
	#10 counter$count = 90713;
	#10 counter$count = 90714;
	#10 counter$count = 90715;
	#10 counter$count = 90716;
	#10 counter$count = 90717;
	#10 counter$count = 90718;
	#10 counter$count = 90719;
	#10 counter$count = 90720;
	#10 counter$count = 90721;
	#10 counter$count = 90722;
	#10 counter$count = 90723;
	#10 counter$count = 90724;
	#10 counter$count = 90725;
	#10 counter$count = 90726;
	#10 counter$count = 90727;
	#10 counter$count = 90728;
	#10 counter$count = 90729;
	#10 counter$count = 90730;
	#10 counter$count = 90731;
	#10 counter$count = 90732;
	#10 counter$count = 90733;
	#10 counter$count = 90734;
	#10 counter$count = 90735;
	#10 counter$count = 90736;
	#10 counter$count = 90737;
	#10 counter$count = 90738;
	#10 counter$count = 90739;
	#10 counter$count = 90740;
	#10 counter$count = 90741;
	#10 counter$count = 90742;
	#10 counter$count = 90743;
	#10 counter$count = 90744;
	#10 counter$count = 90745;
	#10 counter$count = 90746;
	#10 counter$count = 90747;
	#10 counter$count = 90748;
	#10 counter$count = 90749;
	#10 counter$count = 90750;
	#10 counter$count = 90751;
	#10 counter$count = 90752;
	#10 counter$count = 90753;
	#10 counter$count = 90754;
	#10 counter$count = 90755;
	#10 counter$count = 90756;
	#10 counter$count = 90757;
	#10 counter$count = 90758;
	#10 counter$count = 90759;
	#10 counter$count = 90760;
	#10 counter$count = 90761;
	#10 counter$count = 90762;
	#10 counter$count = 90763;
	#10 counter$count = 90764;
	#10 counter$count = 90765;
	#10 counter$count = 90766;
	#10 counter$count = 90767;
	#10 counter$count = 90768;
	#10 counter$count = 90769;
	#10 counter$count = 90770;
	#10 counter$count = 90771;
	#10 counter$count = 90772;
	#10 counter$count = 90773;
	#10 counter$count = 90774;
	#10 counter$count = 90775;
	#10 counter$count = 90776;
	#10 counter$count = 90777;
	#10 counter$count = 90778;
	#10 counter$count = 90779;
	#10 counter$count = 90780;
	#10 counter$count = 90781;
	#10 counter$count = 90782;
	#10 counter$count = 90783;
	#10 counter$count = 90784;
	#10 counter$count = 90785;
	#10 counter$count = 90786;
	#10 counter$count = 90787;
	#10 counter$count = 90788;
	#10 counter$count = 90789;
	#10 counter$count = 90790;
	#10 counter$count = 90791;
	#10 counter$count = 90792;
	#10 counter$count = 90793;
	#10 counter$count = 90794;
	#10 counter$count = 90795;
	#10 counter$count = 90796;
	#10 counter$count = 90797;
	#10 counter$count = 90798;
	#10 counter$count = 90799;
	#10 counter$count = 90800;
	#10 counter$count = 90801;
	#10 counter$count = 90802;
	#10 counter$count = 90803;
	#10 counter$count = 90804;
	#10 counter$count = 90805;
	#10 counter$count = 90806;
	#10 counter$count = 90807;
	#10 counter$count = 90808;
	#10 counter$count = 90809;
	#10 counter$count = 90810;
	#10 counter$count = 90811;
	#10 counter$count = 90812;
	#10 counter$count = 90813;
	#10 counter$count = 90814;
	#10 counter$count = 90815;
	#10 counter$count = 90816;
	#10 counter$count = 90817;
	#10 counter$count = 90818;
	#10 counter$count = 90819;
	#10 counter$count = 90820;
	#10 counter$count = 90821;
	#10 counter$count = 90822;
	#10 counter$count = 90823;
	#10 counter$count = 90824;
	#10 counter$count = 90825;
	#10 counter$count = 90826;
	#10 counter$count = 90827;
	#10 counter$count = 90828;
	#10 counter$count = 90829;
	#10 counter$count = 90830;
	#10 counter$count = 90831;
	#10 counter$count = 90832;
	#10 counter$count = 90833;
	#10 counter$count = 90834;
	#10 counter$count = 90835;
	#10 counter$count = 90836;
	#10 counter$count = 90837;
	#10 counter$count = 90838;
	#10 counter$count = 90839;
	#10 counter$count = 90840;
	#10 counter$count = 90841;
	#10 counter$count = 90842;
	#10 counter$count = 90843;
	#10 counter$count = 90844;
	#10 counter$count = 90845;
	#10 counter$count = 90846;
	#10 counter$count = 90847;
	#10 counter$count = 90848;
	#10 counter$count = 90849;
	#10 counter$count = 90850;
	#10 counter$count = 90851;
	#10 counter$count = 90852;
	#10 counter$count = 90853;
	#10 counter$count = 90854;
	#10 counter$count = 90855;
	#10 counter$count = 90856;
	#10 counter$count = 90857;
	#10 counter$count = 90858;
	#10 counter$count = 90859;
	#10 counter$count = 90860;
	#10 counter$count = 90861;
	#10 counter$count = 90862;
	#10 counter$count = 90863;
	#10 counter$count = 90864;
	#10 counter$count = 90865;
	#10 counter$count = 90866;
	#10 counter$count = 90867;
	#10 counter$count = 90868;
	#10 counter$count = 90869;
	#10 counter$count = 90870;
	#10 counter$count = 90871;
	#10 counter$count = 90872;
	#10 counter$count = 90873;
	#10 counter$count = 90874;
	#10 counter$count = 90875;
	#10 counter$count = 90876;
	#10 counter$count = 90877;
	#10 counter$count = 90878;
	#10 counter$count = 90879;
	#10 counter$count = 90880;
	#10 counter$count = 90881;
	#10 counter$count = 90882;
	#10 counter$count = 90883;
	#10 counter$count = 90884;
	#10 counter$count = 90885;
	#10 counter$count = 90886;
	#10 counter$count = 90887;
	#10 counter$count = 90888;
	#10 counter$count = 90889;
	#10 counter$count = 90890;
	#10 counter$count = 90891;
	#10 counter$count = 90892;
	#10 counter$count = 90893;
	#10 counter$count = 90894;
	#10 counter$count = 90895;
	#10 counter$count = 90896;
	#10 counter$count = 90897;
	#10 counter$count = 90898;
	#10 counter$count = 90899;
	#10 counter$count = 90900;
	#10 counter$count = 90901;
	#10 counter$count = 90902;
	#10 counter$count = 90903;
	#10 counter$count = 90904;
	#10 counter$count = 90905;
	#10 counter$count = 90906;
	#10 counter$count = 90907;
	#10 counter$count = 90908;
	#10 counter$count = 90909;
	#10 counter$count = 90910;
	#10 counter$count = 90911;
	#10 counter$count = 90912;
	#10 counter$count = 90913;
	#10 counter$count = 90914;
	#10 counter$count = 90915;
	#10 counter$count = 90916;
	#10 counter$count = 90917;
	#10 counter$count = 90918;
	#10 counter$count = 90919;
	#10 counter$count = 90920;
	#10 counter$count = 90921;
	#10 counter$count = 90922;
	#10 counter$count = 90923;
	#10 counter$count = 90924;
	#10 counter$count = 90925;
	#10 counter$count = 90926;
	#10 counter$count = 90927;
	#10 counter$count = 90928;
	#10 counter$count = 90929;
	#10 counter$count = 90930;
	#10 counter$count = 90931;
	#10 counter$count = 90932;
	#10 counter$count = 90933;
	#10 counter$count = 90934;
	#10 counter$count = 90935;
	#10 counter$count = 90936;
	#10 counter$count = 90937;
	#10 counter$count = 90938;
	#10 counter$count = 90939;
	#10 counter$count = 90940;
	#10 counter$count = 90941;
	#10 counter$count = 90942;
	#10 counter$count = 90943;
	#10 counter$count = 90944;
	#10 counter$count = 90945;
	#10 counter$count = 90946;
	#10 counter$count = 90947;
	#10 counter$count = 90948;
	#10 counter$count = 90949;
	#10 counter$count = 90950;
	#10 counter$count = 90951;
	#10 counter$count = 90952;
	#10 counter$count = 90953;
	#10 counter$count = 90954;
	#10 counter$count = 90955;
	#10 counter$count = 90956;
	#10 counter$count = 90957;
	#10 counter$count = 90958;
	#10 counter$count = 90959;
	#10 counter$count = 90960;
	#10 counter$count = 90961;
	#10 counter$count = 90962;
	#10 counter$count = 90963;
	#10 counter$count = 90964;
	#10 counter$count = 90965;
	#10 counter$count = 90966;
	#10 counter$count = 90967;
	#10 counter$count = 90968;
	#10 counter$count = 90969;
	#10 counter$count = 90970;
	#10 counter$count = 90971;
	#10 counter$count = 90972;
	#10 counter$count = 90973;
	#10 counter$count = 90974;
	#10 counter$count = 90975;
	#10 counter$count = 90976;
	#10 counter$count = 90977;
	#10 counter$count = 90978;
	#10 counter$count = 90979;
	#10 counter$count = 90980;
	#10 counter$count = 90981;
	#10 counter$count = 90982;
	#10 counter$count = 90983;
	#10 counter$count = 90984;
	#10 counter$count = 90985;
	#10 counter$count = 90986;
	#10 counter$count = 90987;
	#10 counter$count = 90988;
	#10 counter$count = 90989;
	#10 counter$count = 90990;
	#10 counter$count = 90991;
	#10 counter$count = 90992;
	#10 counter$count = 90993;
	#10 counter$count = 90994;
	#10 counter$count = 90995;
	#10 counter$count = 90996;
	#10 counter$count = 90997;
	#10 counter$count = 90998;
	#10 counter$count = 90999;
	#10 counter$count = 91000;
	#10 counter$count = 91001;
	#10 counter$count = 91002;
	#10 counter$count = 91003;
	#10 counter$count = 91004;
	#10 counter$count = 91005;
	#10 counter$count = 91006;
	#10 counter$count = 91007;
	#10 counter$count = 91008;
	#10 counter$count = 91009;
	#10 counter$count = 91010;
	#10 counter$count = 91011;
	#10 counter$count = 91012;
	#10 counter$count = 91013;
	#10 counter$count = 91014;
	#10 counter$count = 91015;
	#10 counter$count = 91016;
	#10 counter$count = 91017;
	#10 counter$count = 91018;
	#10 counter$count = 91019;
	#10 counter$count = 91020;
	#10 counter$count = 91021;
	#10 counter$count = 91022;
	#10 counter$count = 91023;
	#10 counter$count = 91024;
	#10 counter$count = 91025;
	#10 counter$count = 91026;
	#10 counter$count = 91027;
	#10 counter$count = 91028;
	#10 counter$count = 91029;
	#10 counter$count = 91030;
	#10 counter$count = 91031;
	#10 counter$count = 91032;
	#10 counter$count = 91033;
	#10 counter$count = 91034;
	#10 counter$count = 91035;
	#10 counter$count = 91036;
	#10 counter$count = 91037;
	#10 counter$count = 91038;
	#10 counter$count = 91039;
	#10 counter$count = 91040;
	#10 counter$count = 91041;
	#10 counter$count = 91042;
	#10 counter$count = 91043;
	#10 counter$count = 91044;
	#10 counter$count = 91045;
	#10 counter$count = 91046;
	#10 counter$count = 91047;
	#10 counter$count = 91048;
	#10 counter$count = 91049;
	#10 counter$count = 91050;
	#10 counter$count = 91051;
	#10 counter$count = 91052;
	#10 counter$count = 91053;
	#10 counter$count = 91054;
	#10 counter$count = 91055;
	#10 counter$count = 91056;
	#10 counter$count = 91057;
	#10 counter$count = 91058;
	#10 counter$count = 91059;
	#10 counter$count = 91060;
	#10 counter$count = 91061;
	#10 counter$count = 91062;
	#10 counter$count = 91063;
	#10 counter$count = 91064;
	#10 counter$count = 91065;
	#10 counter$count = 91066;
	#10 counter$count = 91067;
	#10 counter$count = 91068;
	#10 counter$count = 91069;
	#10 counter$count = 91070;
	#10 counter$count = 91071;
	#10 counter$count = 91072;
	#10 counter$count = 91073;
	#10 counter$count = 91074;
	#10 counter$count = 91075;
	#10 counter$count = 91076;
	#10 counter$count = 91077;
	#10 counter$count = 91078;
	#10 counter$count = 91079;
	#10 counter$count = 91080;
	#10 counter$count = 91081;
	#10 counter$count = 91082;
	#10 counter$count = 91083;
	#10 counter$count = 91084;
	#10 counter$count = 91085;
	#10 counter$count = 91086;
	#10 counter$count = 91087;
	#10 counter$count = 91088;
	#10 counter$count = 91089;
	#10 counter$count = 91090;
	#10 counter$count = 91091;
	#10 counter$count = 91092;
	#10 counter$count = 91093;
	#10 counter$count = 91094;
	#10 counter$count = 91095;
	#10 counter$count = 91096;
	#10 counter$count = 91097;
	#10 counter$count = 91098;
	#10 counter$count = 91099;
	#10 counter$count = 91100;
	#10 counter$count = 91101;
	#10 counter$count = 91102;
	#10 counter$count = 91103;
	#10 counter$count = 91104;
	#10 counter$count = 91105;
	#10 counter$count = 91106;
	#10 counter$count = 91107;
	#10 counter$count = 91108;
	#10 counter$count = 91109;
	#10 counter$count = 91110;
	#10 counter$count = 91111;
	#10 counter$count = 91112;
	#10 counter$count = 91113;
	#10 counter$count = 91114;
	#10 counter$count = 91115;
	#10 counter$count = 91116;
	#10 counter$count = 91117;
	#10 counter$count = 91118;
	#10 counter$count = 91119;
	#10 counter$count = 91120;
	#10 counter$count = 91121;
	#10 counter$count = 91122;
	#10 counter$count = 91123;
	#10 counter$count = 91124;
	#10 counter$count = 91125;
	#10 counter$count = 91126;
	#10 counter$count = 91127;
	#10 counter$count = 91128;
	#10 counter$count = 91129;
	#10 counter$count = 91130;
	#10 counter$count = 91131;
	#10 counter$count = 91132;
	#10 counter$count = 91133;
	#10 counter$count = 91134;
	#10 counter$count = 91135;
	#10 counter$count = 91136;
	#10 counter$count = 91137;
	#10 counter$count = 91138;
	#10 counter$count = 91139;
	#10 counter$count = 91140;
	#10 counter$count = 91141;
	#10 counter$count = 91142;
	#10 counter$count = 91143;
	#10 counter$count = 91144;
	#10 counter$count = 91145;
	#10 counter$count = 91146;
	#10 counter$count = 91147;
	#10 counter$count = 91148;
	#10 counter$count = 91149;
	#10 counter$count = 91150;
	#10 counter$count = 91151;
	#10 counter$count = 91152;
	#10 counter$count = 91153;
	#10 counter$count = 91154;
	#10 counter$count = 91155;
	#10 counter$count = 91156;
	#10 counter$count = 91157;
	#10 counter$count = 91158;
	#10 counter$count = 91159;
	#10 counter$count = 91160;
	#10 counter$count = 91161;
	#10 counter$count = 91162;
	#10 counter$count = 91163;
	#10 counter$count = 91164;
	#10 counter$count = 91165;
	#10 counter$count = 91166;
	#10 counter$count = 91167;
	#10 counter$count = 91168;
	#10 counter$count = 91169;
	#10 counter$count = 91170;
	#10 counter$count = 91171;
	#10 counter$count = 91172;
	#10 counter$count = 91173;
	#10 counter$count = 91174;
	#10 counter$count = 91175;
	#10 counter$count = 91176;
	#10 counter$count = 91177;
	#10 counter$count = 91178;
	#10 counter$count = 91179;
	#10 counter$count = 91180;
	#10 counter$count = 91181;
	#10 counter$count = 91182;
	#10 counter$count = 91183;
	#10 counter$count = 91184;
	#10 counter$count = 91185;
	#10 counter$count = 91186;
	#10 counter$count = 91187;
	#10 counter$count = 91188;
	#10 counter$count = 91189;
	#10 counter$count = 91190;
	#10 counter$count = 91191;
	#10 counter$count = 91192;
	#10 counter$count = 91193;
	#10 counter$count = 91194;
	#10 counter$count = 91195;
	#10 counter$count = 91196;
	#10 counter$count = 91197;
	#10 counter$count = 91198;
	#10 counter$count = 91199;
	#10 counter$count = 91200;
	#10 counter$count = 91201;
	#10 counter$count = 91202;
	#10 counter$count = 91203;
	#10 counter$count = 91204;
	#10 counter$count = 91205;
	#10 counter$count = 91206;
	#10 counter$count = 91207;
	#10 counter$count = 91208;
	#10 counter$count = 91209;
	#10 counter$count = 91210;
	#10 counter$count = 91211;
	#10 counter$count = 91212;
	#10 counter$count = 91213;
	#10 counter$count = 91214;
	#10 counter$count = 91215;
	#10 counter$count = 91216;
	#10 counter$count = 91217;
	#10 counter$count = 91218;
	#10 counter$count = 91219;
	#10 counter$count = 91220;
	#10 counter$count = 91221;
	#10 counter$count = 91222;
	#10 counter$count = 91223;
	#10 counter$count = 91224;
	#10 counter$count = 91225;
	#10 counter$count = 91226;
	#10 counter$count = 91227;
	#10 counter$count = 91228;
	#10 counter$count = 91229;
	#10 counter$count = 91230;
	#10 counter$count = 91231;
	#10 counter$count = 91232;
	#10 counter$count = 91233;
	#10 counter$count = 91234;
	#10 counter$count = 91235;
	#10 counter$count = 91236;
	#10 counter$count = 91237;
	#10 counter$count = 91238;
	#10 counter$count = 91239;
	#10 counter$count = 91240;
	#10 counter$count = 91241;
	#10 counter$count = 91242;
	#10 counter$count = 91243;
	#10 counter$count = 91244;
	#10 counter$count = 91245;
	#10 counter$count = 91246;
	#10 counter$count = 91247;
	#10 counter$count = 91248;
	#10 counter$count = 91249;
	#10 counter$count = 91250;
	#10 counter$count = 91251;
	#10 counter$count = 91252;
	#10 counter$count = 91253;
	#10 counter$count = 91254;
	#10 counter$count = 91255;
	#10 counter$count = 91256;
	#10 counter$count = 91257;
	#10 counter$count = 91258;
	#10 counter$count = 91259;
	#10 counter$count = 91260;
	#10 counter$count = 91261;
	#10 counter$count = 91262;
	#10 counter$count = 91263;
	#10 counter$count = 91264;
	#10 counter$count = 91265;
	#10 counter$count = 91266;
	#10 counter$count = 91267;
	#10 counter$count = 91268;
	#10 counter$count = 91269;
	#10 counter$count = 91270;
	#10 counter$count = 91271;
	#10 counter$count = 91272;
	#10 counter$count = 91273;
	#10 counter$count = 91274;
	#10 counter$count = 91275;
	#10 counter$count = 91276;
	#10 counter$count = 91277;
	#10 counter$count = 91278;
	#10 counter$count = 91279;
	#10 counter$count = 91280;
	#10 counter$count = 91281;
	#10 counter$count = 91282;
	#10 counter$count = 91283;
	#10 counter$count = 91284;
	#10 counter$count = 91285;
	#10 counter$count = 91286;
	#10 counter$count = 91287;
	#10 counter$count = 91288;
	#10 counter$count = 91289;
	#10 counter$count = 91290;
	#10 counter$count = 91291;
	#10 counter$count = 91292;
	#10 counter$count = 91293;
	#10 counter$count = 91294;
	#10 counter$count = 91295;
	#10 counter$count = 91296;
	#10 counter$count = 91297;
	#10 counter$count = 91298;
	#10 counter$count = 91299;
	#10 counter$count = 91300;
	#10 counter$count = 91301;
	#10 counter$count = 91302;
	#10 counter$count = 91303;
	#10 counter$count = 91304;
	#10 counter$count = 91305;
	#10 counter$count = 91306;
	#10 counter$count = 91307;
	#10 counter$count = 91308;
	#10 counter$count = 91309;
	#10 counter$count = 91310;
	#10 counter$count = 91311;
	#10 counter$count = 91312;
	#10 counter$count = 91313;
	#10 counter$count = 91314;
	#10 counter$count = 91315;
	#10 counter$count = 91316;
	#10 counter$count = 91317;
	#10 counter$count = 91318;
	#10 counter$count = 91319;
	#10 counter$count = 91320;
	#10 counter$count = 91321;
	#10 counter$count = 91322;
	#10 counter$count = 91323;
	#10 counter$count = 91324;
	#10 counter$count = 91325;
	#10 counter$count = 91326;
	#10 counter$count = 91327;
	#10 counter$count = 91328;
	#10 counter$count = 91329;
	#10 counter$count = 91330;
	#10 counter$count = 91331;
	#10 counter$count = 91332;
	#10 counter$count = 91333;
	#10 counter$count = 91334;
	#10 counter$count = 91335;
	#10 counter$count = 91336;
	#10 counter$count = 91337;
	#10 counter$count = 91338;
	#10 counter$count = 91339;
	#10 counter$count = 91340;
	#10 counter$count = 91341;
	#10 counter$count = 91342;
	#10 counter$count = 91343;
	#10 counter$count = 91344;
	#10 counter$count = 91345;
	#10 counter$count = 91346;
	#10 counter$count = 91347;
	#10 counter$count = 91348;
	#10 counter$count = 91349;
	#10 counter$count = 91350;
	#10 counter$count = 91351;
	#10 counter$count = 91352;
	#10 counter$count = 91353;
	#10 counter$count = 91354;
	#10 counter$count = 91355;
	#10 counter$count = 91356;
	#10 counter$count = 91357;
	#10 counter$count = 91358;
	#10 counter$count = 91359;
	#10 counter$count = 91360;
	#10 counter$count = 91361;
	#10 counter$count = 91362;
	#10 counter$count = 91363;
	#10 counter$count = 91364;
	#10 counter$count = 91365;
	#10 counter$count = 91366;
	#10 counter$count = 91367;
	#10 counter$count = 91368;
	#10 counter$count = 91369;
	#10 counter$count = 91370;
	#10 counter$count = 91371;
	#10 counter$count = 91372;
	#10 counter$count = 91373;
	#10 counter$count = 91374;
	#10 counter$count = 91375;
	#10 counter$count = 91376;
	#10 counter$count = 91377;
	#10 counter$count = 91378;
	#10 counter$count = 91379;
	#10 counter$count = 91380;
	#10 counter$count = 91381;
	#10 counter$count = 91382;
	#10 counter$count = 91383;
	#10 counter$count = 91384;
	#10 counter$count = 91385;
	#10 counter$count = 91386;
	#10 counter$count = 91387;
	#10 counter$count = 91388;
	#10 counter$count = 91389;
	#10 counter$count = 91390;
	#10 counter$count = 91391;
	#10 counter$count = 91392;
	#10 counter$count = 91393;
	#10 counter$count = 91394;
	#10 counter$count = 91395;
	#10 counter$count = 91396;
	#10 counter$count = 91397;
	#10 counter$count = 91398;
	#10 counter$count = 91399;
	#10 counter$count = 91400;
	#10 counter$count = 91401;
	#10 counter$count = 91402;
	#10 counter$count = 91403;
	#10 counter$count = 91404;
	#10 counter$count = 91405;
	#10 counter$count = 91406;
	#10 counter$count = 91407;
	#10 counter$count = 91408;
	#10 counter$count = 91409;
	#10 counter$count = 91410;
	#10 counter$count = 91411;
	#10 counter$count = 91412;
	#10 counter$count = 91413;
	#10 counter$count = 91414;
	#10 counter$count = 91415;
	#10 counter$count = 91416;
	#10 counter$count = 91417;
	#10 counter$count = 91418;
	#10 counter$count = 91419;
	#10 counter$count = 91420;
	#10 counter$count = 91421;
	#10 counter$count = 91422;
	#10 counter$count = 91423;
	#10 counter$count = 91424;
	#10 counter$count = 91425;
	#10 counter$count = 91426;
	#10 counter$count = 91427;
	#10 counter$count = 91428;
	#10 counter$count = 91429;
	#10 counter$count = 91430;
	#10 counter$count = 91431;
	#10 counter$count = 91432;
	#10 counter$count = 91433;
	#10 counter$count = 91434;
	#10 counter$count = 91435;
	#10 counter$count = 91436;
	#10 counter$count = 91437;
	#10 counter$count = 91438;
	#10 counter$count = 91439;
	#10 counter$count = 91440;
	#10 counter$count = 91441;
	#10 counter$count = 91442;
	#10 counter$count = 91443;
	#10 counter$count = 91444;
	#10 counter$count = 91445;
	#10 counter$count = 91446;
	#10 counter$count = 91447;
	#10 counter$count = 91448;
	#10 counter$count = 91449;
	#10 counter$count = 91450;
	#10 counter$count = 91451;
	#10 counter$count = 91452;
	#10 counter$count = 91453;
	#10 counter$count = 91454;
	#10 counter$count = 91455;
	#10 counter$count = 91456;
	#10 counter$count = 91457;
	#10 counter$count = 91458;
	#10 counter$count = 91459;
	#10 counter$count = 91460;
	#10 counter$count = 91461;
	#10 counter$count = 91462;
	#10 counter$count = 91463;
	#10 counter$count = 91464;
	#10 counter$count = 91465;
	#10 counter$count = 91466;
	#10 counter$count = 91467;
	#10 counter$count = 91468;
	#10 counter$count = 91469;
	#10 counter$count = 91470;
	#10 counter$count = 91471;
	#10 counter$count = 91472;
	#10 counter$count = 91473;
	#10 counter$count = 91474;
	#10 counter$count = 91475;
	#10 counter$count = 91476;
	#10 counter$count = 91477;
	#10 counter$count = 91478;
	#10 counter$count = 91479;
	#10 counter$count = 91480;
	#10 counter$count = 91481;
	#10 counter$count = 91482;
	#10 counter$count = 91483;
	#10 counter$count = 91484;
	#10 counter$count = 91485;
	#10 counter$count = 91486;
	#10 counter$count = 91487;
	#10 counter$count = 91488;
	#10 counter$count = 91489;
	#10 counter$count = 91490;
	#10 counter$count = 91491;
	#10 counter$count = 91492;
	#10 counter$count = 91493;
	#10 counter$count = 91494;
	#10 counter$count = 91495;
	#10 counter$count = 91496;
	#10 counter$count = 91497;
	#10 counter$count = 91498;
	#10 counter$count = 91499;
	#10 counter$count = 91500;
	#10 counter$count = 91501;
	#10 counter$count = 91502;
	#10 counter$count = 91503;
	#10 counter$count = 91504;
	#10 counter$count = 91505;
	#10 counter$count = 91506;
	#10 counter$count = 91507;
	#10 counter$count = 91508;
	#10 counter$count = 91509;
	#10 counter$count = 91510;
	#10 counter$count = 91511;
	#10 counter$count = 91512;
	#10 counter$count = 91513;
	#10 counter$count = 91514;
	#10 counter$count = 91515;
	#10 counter$count = 91516;
	#10 counter$count = 91517;
	#10 counter$count = 91518;
	#10 counter$count = 91519;
	#10 counter$count = 91520;
	#10 counter$count = 91521;
	#10 counter$count = 91522;
	#10 counter$count = 91523;
	#10 counter$count = 91524;
	#10 counter$count = 91525;
	#10 counter$count = 91526;
	#10 counter$count = 91527;
	#10 counter$count = 91528;
	#10 counter$count = 91529;
	#10 counter$count = 91530;
	#10 counter$count = 91531;
	#10 counter$count = 91532;
	#10 counter$count = 91533;
	#10 counter$count = 91534;
	#10 counter$count = 91535;
	#10 counter$count = 91536;
	#10 counter$count = 91537;
	#10 counter$count = 91538;
	#10 counter$count = 91539;
	#10 counter$count = 91540;
	#10 counter$count = 91541;
	#10 counter$count = 91542;
	#10 counter$count = 91543;
	#10 counter$count = 91544;
	#10 counter$count = 91545;
	#10 counter$count = 91546;
	#10 counter$count = 91547;
	#10 counter$count = 91548;
	#10 counter$count = 91549;
	#10 counter$count = 91550;
	#10 counter$count = 91551;
	#10 counter$count = 91552;
	#10 counter$count = 91553;
	#10 counter$count = 91554;
	#10 counter$count = 91555;
	#10 counter$count = 91556;
	#10 counter$count = 91557;
	#10 counter$count = 91558;
	#10 counter$count = 91559;
	#10 counter$count = 91560;
	#10 counter$count = 91561;
	#10 counter$count = 91562;
	#10 counter$count = 91563;
	#10 counter$count = 91564;
	#10 counter$count = 91565;
	#10 counter$count = 91566;
	#10 counter$count = 91567;
	#10 counter$count = 91568;
	#10 counter$count = 91569;
	#10 counter$count = 91570;
	#10 counter$count = 91571;
	#10 counter$count = 91572;
	#10 counter$count = 91573;
	#10 counter$count = 91574;
	#10 counter$count = 91575;
	#10 counter$count = 91576;
	#10 counter$count = 91577;
	#10 counter$count = 91578;
	#10 counter$count = 91579;
	#10 counter$count = 91580;
	#10 counter$count = 91581;
	#10 counter$count = 91582;
	#10 counter$count = 91583;
	#10 counter$count = 91584;
	#10 counter$count = 91585;
	#10 counter$count = 91586;
	#10 counter$count = 91587;
	#10 counter$count = 91588;
	#10 counter$count = 91589;
	#10 counter$count = 91590;
	#10 counter$count = 91591;
	#10 counter$count = 91592;
	#10 counter$count = 91593;
	#10 counter$count = 91594;
	#10 counter$count = 91595;
	#10 counter$count = 91596;
	#10 counter$count = 91597;
	#10 counter$count = 91598;
	#10 counter$count = 91599;
	#10 counter$count = 91600;
	#10 counter$count = 91601;
	#10 counter$count = 91602;
	#10 counter$count = 91603;
	#10 counter$count = 91604;
	#10 counter$count = 91605;
	#10 counter$count = 91606;
	#10 counter$count = 91607;
	#10 counter$count = 91608;
	#10 counter$count = 91609;
	#10 counter$count = 91610;
	#10 counter$count = 91611;
	#10 counter$count = 91612;
	#10 counter$count = 91613;
	#10 counter$count = 91614;
	#10 counter$count = 91615;
	#10 counter$count = 91616;
	#10 counter$count = 91617;
	#10 counter$count = 91618;
	#10 counter$count = 91619;
	#10 counter$count = 91620;
	#10 counter$count = 91621;
	#10 counter$count = 91622;
	#10 counter$count = 91623;
	#10 counter$count = 91624;
	#10 counter$count = 91625;
	#10 counter$count = 91626;
	#10 counter$count = 91627;
	#10 counter$count = 91628;
	#10 counter$count = 91629;
	#10 counter$count = 91630;
	#10 counter$count = 91631;
	#10 counter$count = 91632;
	#10 counter$count = 91633;
	#10 counter$count = 91634;
	#10 counter$count = 91635;
	#10 counter$count = 91636;
	#10 counter$count = 91637;
	#10 counter$count = 91638;
	#10 counter$count = 91639;
	#10 counter$count = 91640;
	#10 counter$count = 91641;
	#10 counter$count = 91642;
	#10 counter$count = 91643;
	#10 counter$count = 91644;
	#10 counter$count = 91645;
	#10 counter$count = 91646;
	#10 counter$count = 91647;
	#10 counter$count = 91648;
	#10 counter$count = 91649;
	#10 counter$count = 91650;
	#10 counter$count = 91651;
	#10 counter$count = 91652;
	#10 counter$count = 91653;
	#10 counter$count = 91654;
	#10 counter$count = 91655;
	#10 counter$count = 91656;
	#10 counter$count = 91657;
	#10 counter$count = 91658;
	#10 counter$count = 91659;
	#10 counter$count = 91660;
	#10 counter$count = 91661;
	#10 counter$count = 91662;
	#10 counter$count = 91663;
	#10 counter$count = 91664;
	#10 counter$count = 91665;
	#10 counter$count = 91666;
	#10 counter$count = 91667;
	#10 counter$count = 91668;
	#10 counter$count = 91669;
	#10 counter$count = 91670;
	#10 counter$count = 91671;
	#10 counter$count = 91672;
	#10 counter$count = 91673;
	#10 counter$count = 91674;
	#10 counter$count = 91675;
	#10 counter$count = 91676;
	#10 counter$count = 91677;
	#10 counter$count = 91678;
	#10 counter$count = 91679;
	#10 counter$count = 91680;
	#10 counter$count = 91681;
	#10 counter$count = 91682;
	#10 counter$count = 91683;
	#10 counter$count = 91684;
	#10 counter$count = 91685;
	#10 counter$count = 91686;
	#10 counter$count = 91687;
	#10 counter$count = 91688;
	#10 counter$count = 91689;
	#10 counter$count = 91690;
	#10 counter$count = 91691;
	#10 counter$count = 91692;
	#10 counter$count = 91693;
	#10 counter$count = 91694;
	#10 counter$count = 91695;
	#10 counter$count = 91696;
	#10 counter$count = 91697;
	#10 counter$count = 91698;
	#10 counter$count = 91699;
	#10 counter$count = 91700;
	#10 counter$count = 91701;
	#10 counter$count = 91702;
	#10 counter$count = 91703;
	#10 counter$count = 91704;
	#10 counter$count = 91705;
	#10 counter$count = 91706;
	#10 counter$count = 91707;
	#10 counter$count = 91708;
	#10 counter$count = 91709;
	#10 counter$count = 91710;
	#10 counter$count = 91711;
	#10 counter$count = 91712;
	#10 counter$count = 91713;
	#10 counter$count = 91714;
	#10 counter$count = 91715;
	#10 counter$count = 91716;
	#10 counter$count = 91717;
	#10 counter$count = 91718;
	#10 counter$count = 91719;
	#10 counter$count = 91720;
	#10 counter$count = 91721;
	#10 counter$count = 91722;
	#10 counter$count = 91723;
	#10 counter$count = 91724;
	#10 counter$count = 91725;
	#10 counter$count = 91726;
	#10 counter$count = 91727;
	#10 counter$count = 91728;
	#10 counter$count = 91729;
	#10 counter$count = 91730;
	#10 counter$count = 91731;
	#10 counter$count = 91732;
	#10 counter$count = 91733;
	#10 counter$count = 91734;
	#10 counter$count = 91735;
	#10 counter$count = 91736;
	#10 counter$count = 91737;
	#10 counter$count = 91738;
	#10 counter$count = 91739;
	#10 counter$count = 91740;
	#10 counter$count = 91741;
	#10 counter$count = 91742;
	#10 counter$count = 91743;
	#10 counter$count = 91744;
	#10 counter$count = 91745;
	#10 counter$count = 91746;
	#10 counter$count = 91747;
	#10 counter$count = 91748;
	#10 counter$count = 91749;
	#10 counter$count = 91750;
	#10 counter$count = 91751;
	#10 counter$count = 91752;
	#10 counter$count = 91753;
	#10 counter$count = 91754;
	#10 counter$count = 91755;
	#10 counter$count = 91756;
	#10 counter$count = 91757;
	#10 counter$count = 91758;
	#10 counter$count = 91759;
	#10 counter$count = 91760;
	#10 counter$count = 91761;
	#10 counter$count = 91762;
	#10 counter$count = 91763;
	#10 counter$count = 91764;
	#10 counter$count = 91765;
	#10 counter$count = 91766;
	#10 counter$count = 91767;
	#10 counter$count = 91768;
	#10 counter$count = 91769;
	#10 counter$count = 91770;
	#10 counter$count = 91771;
	#10 counter$count = 91772;
	#10 counter$count = 91773;
	#10 counter$count = 91774;
	#10 counter$count = 91775;
	#10 counter$count = 91776;
	#10 counter$count = 91777;
	#10 counter$count = 91778;
	#10 counter$count = 91779;
	#10 counter$count = 91780;
	#10 counter$count = 91781;
	#10 counter$count = 91782;
	#10 counter$count = 91783;
	#10 counter$count = 91784;
	#10 counter$count = 91785;
	#10 counter$count = 91786;
	#10 counter$count = 91787;
	#10 counter$count = 91788;
	#10 counter$count = 91789;
	#10 counter$count = 91790;
	#10 counter$count = 91791;
	#10 counter$count = 91792;
	#10 counter$count = 91793;
	#10 counter$count = 91794;
	#10 counter$count = 91795;
	#10 counter$count = 91796;
	#10 counter$count = 91797;
	#10 counter$count = 91798;
	#10 counter$count = 91799;
	#10 counter$count = 91800;
	#10 counter$count = 91801;
	#10 counter$count = 91802;
	#10 counter$count = 91803;
	#10 counter$count = 91804;
	#10 counter$count = 91805;
	#10 counter$count = 91806;
	#10 counter$count = 91807;
	#10 counter$count = 91808;
	#10 counter$count = 91809;
	#10 counter$count = 91810;
	#10 counter$count = 91811;
	#10 counter$count = 91812;
	#10 counter$count = 91813;
	#10 counter$count = 91814;
	#10 counter$count = 91815;
	#10 counter$count = 91816;
	#10 counter$count = 91817;
	#10 counter$count = 91818;
	#10 counter$count = 91819;
	#10 counter$count = 91820;
	#10 counter$count = 91821;
	#10 counter$count = 91822;
	#10 counter$count = 91823;
	#10 counter$count = 91824;
	#10 counter$count = 91825;
	#10 counter$count = 91826;
	#10 counter$count = 91827;
	#10 counter$count = 91828;
	#10 counter$count = 91829;
	#10 counter$count = 91830;
	#10 counter$count = 91831;
	#10 counter$count = 91832;
	#10 counter$count = 91833;
	#10 counter$count = 91834;
	#10 counter$count = 91835;
	#10 counter$count = 91836;
	#10 counter$count = 91837;
	#10 counter$count = 91838;
	#10 counter$count = 91839;
	#10 counter$count = 91840;
	#10 counter$count = 91841;
	#10 counter$count = 91842;
	#10 counter$count = 91843;
	#10 counter$count = 91844;
	#10 counter$count = 91845;
	#10 counter$count = 91846;
	#10 counter$count = 91847;
	#10 counter$count = 91848;
	#10 counter$count = 91849;
	#10 counter$count = 91850;
	#10 counter$count = 91851;
	#10 counter$count = 91852;
	#10 counter$count = 91853;
	#10 counter$count = 91854;
	#10 counter$count = 91855;
	#10 counter$count = 91856;
	#10 counter$count = 91857;
	#10 counter$count = 91858;
	#10 counter$count = 91859;
	#10 counter$count = 91860;
	#10 counter$count = 91861;
	#10 counter$count = 91862;
	#10 counter$count = 91863;
	#10 counter$count = 91864;
	#10 counter$count = 91865;
	#10 counter$count = 91866;
	#10 counter$count = 91867;
	#10 counter$count = 91868;
	#10 counter$count = 91869;
	#10 counter$count = 91870;
	#10 counter$count = 91871;
	#10 counter$count = 91872;
	#10 counter$count = 91873;
	#10 counter$count = 91874;
	#10 counter$count = 91875;
	#10 counter$count = 91876;
	#10 counter$count = 91877;
	#10 counter$count = 91878;
	#10 counter$count = 91879;
	#10 counter$count = 91880;
	#10 counter$count = 91881;
	#10 counter$count = 91882;
	#10 counter$count = 91883;
	#10 counter$count = 91884;
	#10 counter$count = 91885;
	#10 counter$count = 91886;
	#10 counter$count = 91887;
	#10 counter$count = 91888;
	#10 counter$count = 91889;
	#10 counter$count = 91890;
	#10 counter$count = 91891;
	#10 counter$count = 91892;
	#10 counter$count = 91893;
	#10 counter$count = 91894;
	#10 counter$count = 91895;
	#10 counter$count = 91896;
	#10 counter$count = 91897;
	#10 counter$count = 91898;
	#10 counter$count = 91899;
	#10 counter$count = 91900;
	#10 counter$count = 91901;
	#10 counter$count = 91902;
	#10 counter$count = 91903;
	#10 counter$count = 91904;
	#10 counter$count = 91905;
	#10 counter$count = 91906;
	#10 counter$count = 91907;
	#10 counter$count = 91908;
	#10 counter$count = 91909;
	#10 counter$count = 91910;
	#10 counter$count = 91911;
	#10 counter$count = 91912;
	#10 counter$count = 91913;
	#10 counter$count = 91914;
	#10 counter$count = 91915;
	#10 counter$count = 91916;
	#10 counter$count = 91917;
	#10 counter$count = 91918;
	#10 counter$count = 91919;
	#10 counter$count = 91920;
	#10 counter$count = 91921;
	#10 counter$count = 91922;
	#10 counter$count = 91923;
	#10 counter$count = 91924;
	#10 counter$count = 91925;
	#10 counter$count = 91926;
	#10 counter$count = 91927;
	#10 counter$count = 91928;
	#10 counter$count = 91929;
	#10 counter$count = 91930;
	#10 counter$count = 91931;
	#10 counter$count = 91932;
	#10 counter$count = 91933;
	#10 counter$count = 91934;
	#10 counter$count = 91935;
	#10 counter$count = 91936;
	#10 counter$count = 91937;
	#10 counter$count = 91938;
	#10 counter$count = 91939;
	#10 counter$count = 91940;
	#10 counter$count = 91941;
	#10 counter$count = 91942;
	#10 counter$count = 91943;
	#10 counter$count = 91944;
	#10 counter$count = 91945;
	#10 counter$count = 91946;
	#10 counter$count = 91947;
	#10 counter$count = 91948;
	#10 counter$count = 91949;
	#10 counter$count = 91950;
	#10 counter$count = 91951;
	#10 counter$count = 91952;
	#10 counter$count = 91953;
	#10 counter$count = 91954;
	#10 counter$count = 91955;
	#10 counter$count = 91956;
	#10 counter$count = 91957;
	#10 counter$count = 91958;
	#10 counter$count = 91959;
	#10 counter$count = 91960;
	#10 counter$count = 91961;
	#10 counter$count = 91962;
	#10 counter$count = 91963;
	#10 counter$count = 91964;
	#10 counter$count = 91965;
	#10 counter$count = 91966;
	#10 counter$count = 91967;
	#10 counter$count = 91968;
	#10 counter$count = 91969;
	#10 counter$count = 91970;
	#10 counter$count = 91971;
	#10 counter$count = 91972;
	#10 counter$count = 91973;
	#10 counter$count = 91974;
	#10 counter$count = 91975;
	#10 counter$count = 91976;
	#10 counter$count = 91977;
	#10 counter$count = 91978;
	#10 counter$count = 91979;
	#10 counter$count = 91980;
	#10 counter$count = 91981;
	#10 counter$count = 91982;
	#10 counter$count = 91983;
	#10 counter$count = 91984;
	#10 counter$count = 91985;
	#10 counter$count = 91986;
	#10 counter$count = 91987;
	#10 counter$count = 91988;
	#10 counter$count = 91989;
	#10 counter$count = 91990;
	#10 counter$count = 91991;
	#10 counter$count = 91992;
	#10 counter$count = 91993;
	#10 counter$count = 91994;
	#10 counter$count = 91995;
	#10 counter$count = 91996;
	#10 counter$count = 91997;
	#10 counter$count = 91998;
	#10 counter$count = 91999;
	#10 counter$count = 92000;
	#10 counter$count = 92001;
	#10 counter$count = 92002;
	#10 counter$count = 92003;
	#10 counter$count = 92004;
	#10 counter$count = 92005;
	#10 counter$count = 92006;
	#10 counter$count = 92007;
	#10 counter$count = 92008;
	#10 counter$count = 92009;
	#10 counter$count = 92010;
	#10 counter$count = 92011;
	#10 counter$count = 92012;
	#10 counter$count = 92013;
	#10 counter$count = 92014;
	#10 counter$count = 92015;
	#10 counter$count = 92016;
	#10 counter$count = 92017;
	#10 counter$count = 92018;
	#10 counter$count = 92019;
	#10 counter$count = 92020;
	#10 counter$count = 92021;
	#10 counter$count = 92022;
	#10 counter$count = 92023;
	#10 counter$count = 92024;
	#10 counter$count = 92025;
	#10 counter$count = 92026;
	#10 counter$count = 92027;
	#10 counter$count = 92028;
	#10 counter$count = 92029;
	#10 counter$count = 92030;
	#10 counter$count = 92031;
	#10 counter$count = 92032;
	#10 counter$count = 92033;
	#10 counter$count = 92034;
	#10 counter$count = 92035;
	#10 counter$count = 92036;
	#10 counter$count = 92037;
	#10 counter$count = 92038;
	#10 counter$count = 92039;
	#10 counter$count = 92040;
	#10 counter$count = 92041;
	#10 counter$count = 92042;
	#10 counter$count = 92043;
	#10 counter$count = 92044;
	#10 counter$count = 92045;
	#10 counter$count = 92046;
	#10 counter$count = 92047;
	#10 counter$count = 92048;
	#10 counter$count = 92049;
	#10 counter$count = 92050;
	#10 counter$count = 92051;
	#10 counter$count = 92052;
	#10 counter$count = 92053;
	#10 counter$count = 92054;
	#10 counter$count = 92055;
	#10 counter$count = 92056;
	#10 counter$count = 92057;
	#10 counter$count = 92058;
	#10 counter$count = 92059;
	#10 counter$count = 92060;
	#10 counter$count = 92061;
	#10 counter$count = 92062;
	#10 counter$count = 92063;
	#10 counter$count = 92064;
	#10 counter$count = 92065;
	#10 counter$count = 92066;
	#10 counter$count = 92067;
	#10 counter$count = 92068;
	#10 counter$count = 92069;
	#10 counter$count = 92070;
	#10 counter$count = 92071;
	#10 counter$count = 92072;
	#10 counter$count = 92073;
	#10 counter$count = 92074;
	#10 counter$count = 92075;
	#10 counter$count = 92076;
	#10 counter$count = 92077;
	#10 counter$count = 92078;
	#10 counter$count = 92079;
	#10 counter$count = 92080;
	#10 counter$count = 92081;
	#10 counter$count = 92082;
	#10 counter$count = 92083;
	#10 counter$count = 92084;
	#10 counter$count = 92085;
	#10 counter$count = 92086;
	#10 counter$count = 92087;
	#10 counter$count = 92088;
	#10 counter$count = 92089;
	#10 counter$count = 92090;
	#10 counter$count = 92091;
	#10 counter$count = 92092;
	#10 counter$count = 92093;
	#10 counter$count = 92094;
	#10 counter$count = 92095;
	#10 counter$count = 92096;
	#10 counter$count = 92097;
	#10 counter$count = 92098;
	#10 counter$count = 92099;
	#10 counter$count = 92100;
	#10 counter$count = 92101;
	#10 counter$count = 92102;
	#10 counter$count = 92103;
	#10 counter$count = 92104;
	#10 counter$count = 92105;
	#10 counter$count = 92106;
	#10 counter$count = 92107;
	#10 counter$count = 92108;
	#10 counter$count = 92109;
	#10 counter$count = 92110;
	#10 counter$count = 92111;
	#10 counter$count = 92112;
	#10 counter$count = 92113;
	#10 counter$count = 92114;
	#10 counter$count = 92115;
	#10 counter$count = 92116;
	#10 counter$count = 92117;
	#10 counter$count = 92118;
	#10 counter$count = 92119;
	#10 counter$count = 92120;
	#10 counter$count = 92121;
	#10 counter$count = 92122;
	#10 counter$count = 92123;
	#10 counter$count = 92124;
	#10 counter$count = 92125;
	#10 counter$count = 92126;
	#10 counter$count = 92127;
	#10 counter$count = 92128;
	#10 counter$count = 92129;
	#10 counter$count = 92130;
	#10 counter$count = 92131;
	#10 counter$count = 92132;
	#10 counter$count = 92133;
	#10 counter$count = 92134;
	#10 counter$count = 92135;
	#10 counter$count = 92136;
	#10 counter$count = 92137;
	#10 counter$count = 92138;
	#10 counter$count = 92139;
	#10 counter$count = 92140;
	#10 counter$count = 92141;
	#10 counter$count = 92142;
	#10 counter$count = 92143;
	#10 counter$count = 92144;
	#10 counter$count = 92145;
	#10 counter$count = 92146;
	#10 counter$count = 92147;
	#10 counter$count = 92148;
	#10 counter$count = 92149;
	#10 counter$count = 92150;
	#10 counter$count = 92151;
	#10 counter$count = 92152;
	#10 counter$count = 92153;
	#10 counter$count = 92154;
	#10 counter$count = 92155;
	#10 counter$count = 92156;
	#10 counter$count = 92157;
	#10 counter$count = 92158;
	#10 counter$count = 92159;
	#10 counter$count = 92160;
	#10 counter$count = 92161;
	#10 counter$count = 92162;
	#10 counter$count = 92163;
	#10 counter$count = 92164;
	#10 counter$count = 92165;
	#10 counter$count = 92166;
	#10 counter$count = 92167;
	#10 counter$count = 92168;
	#10 counter$count = 92169;
	#10 counter$count = 92170;
	#10 counter$count = 92171;
	#10 counter$count = 92172;
	#10 counter$count = 92173;
	#10 counter$count = 92174;
	#10 counter$count = 92175;
	#10 counter$count = 92176;
	#10 counter$count = 92177;
	#10 counter$count = 92178;
	#10 counter$count = 92179;
	#10 counter$count = 92180;
	#10 counter$count = 92181;
	#10 counter$count = 92182;
	#10 counter$count = 92183;
	#10 counter$count = 92184;
	#10 counter$count = 92185;
	#10 counter$count = 92186;
	#10 counter$count = 92187;
	#10 counter$count = 92188;
	#10 counter$count = 92189;
	#10 counter$count = 92190;
	#10 counter$count = 92191;
	#10 counter$count = 92192;
	#10 counter$count = 92193;
	#10 counter$count = 92194;
	#10 counter$count = 92195;
	#10 counter$count = 92196;
	#10 counter$count = 92197;
	#10 counter$count = 92198;
	#10 counter$count = 92199;
	#10 counter$count = 92200;
	#10 counter$count = 92201;
	#10 counter$count = 92202;
	#10 counter$count = 92203;
	#10 counter$count = 92204;
	#10 counter$count = 92205;
	#10 counter$count = 92206;
	#10 counter$count = 92207;
	#10 counter$count = 92208;
	#10 counter$count = 92209;
	#10 counter$count = 92210;
	#10 counter$count = 92211;
	#10 counter$count = 92212;
	#10 counter$count = 92213;
	#10 counter$count = 92214;
	#10 counter$count = 92215;
	#10 counter$count = 92216;
	#10 counter$count = 92217;
	#10 counter$count = 92218;
	#10 counter$count = 92219;
	#10 counter$count = 92220;
	#10 counter$count = 92221;
	#10 counter$count = 92222;
	#10 counter$count = 92223;
	#10 counter$count = 92224;
	#10 counter$count = 92225;
	#10 counter$count = 92226;
	#10 counter$count = 92227;
	#10 counter$count = 92228;
	#10 counter$count = 92229;
	#10 counter$count = 92230;
	#10 counter$count = 92231;
	#10 counter$count = 92232;
	#10 counter$count = 92233;
	#10 counter$count = 92234;
	#10 counter$count = 92235;
	#10 counter$count = 92236;
	#10 counter$count = 92237;
	#10 counter$count = 92238;
	#10 counter$count = 92239;
	#10 counter$count = 92240;
	#10 counter$count = 92241;
	#10 counter$count = 92242;
	#10 counter$count = 92243;
	#10 counter$count = 92244;
	#10 counter$count = 92245;
	#10 counter$count = 92246;
	#10 counter$count = 92247;
	#10 counter$count = 92248;
	#10 counter$count = 92249;
	#10 counter$count = 92250;
	#10 counter$count = 92251;
	#10 counter$count = 92252;
	#10 counter$count = 92253;
	#10 counter$count = 92254;
	#10 counter$count = 92255;
	#10 counter$count = 92256;
	#10 counter$count = 92257;
	#10 counter$count = 92258;
	#10 counter$count = 92259;
	#10 counter$count = 92260;
	#10 counter$count = 92261;
	#10 counter$count = 92262;
	#10 counter$count = 92263;
	#10 counter$count = 92264;
	#10 counter$count = 92265;
	#10 counter$count = 92266;
	#10 counter$count = 92267;
	#10 counter$count = 92268;
	#10 counter$count = 92269;
	#10 counter$count = 92270;
	#10 counter$count = 92271;
	#10 counter$count = 92272;
	#10 counter$count = 92273;
	#10 counter$count = 92274;
	#10 counter$count = 92275;
	#10 counter$count = 92276;
	#10 counter$count = 92277;
	#10 counter$count = 92278;
	#10 counter$count = 92279;
	#10 counter$count = 92280;
	#10 counter$count = 92281;
	#10 counter$count = 92282;
	#10 counter$count = 92283;
	#10 counter$count = 92284;
	#10 counter$count = 92285;
	#10 counter$count = 92286;
	#10 counter$count = 92287;
	#10 counter$count = 92288;
	#10 counter$count = 92289;
	#10 counter$count = 92290;
	#10 counter$count = 92291;
	#10 counter$count = 92292;
	#10 counter$count = 92293;
	#10 counter$count = 92294;
	#10 counter$count = 92295;
	#10 counter$count = 92296;
	#10 counter$count = 92297;
	#10 counter$count = 92298;
	#10 counter$count = 92299;
	#10 counter$count = 92300;
	#10 counter$count = 92301;
	#10 counter$count = 92302;
	#10 counter$count = 92303;
	#10 counter$count = 92304;
	#10 counter$count = 92305;
	#10 counter$count = 92306;
	#10 counter$count = 92307;
	#10 counter$count = 92308;
	#10 counter$count = 92309;
	#10 counter$count = 92310;
	#10 counter$count = 92311;
	#10 counter$count = 92312;
	#10 counter$count = 92313;
	#10 counter$count = 92314;
	#10 counter$count = 92315;
	#10 counter$count = 92316;
	#10 counter$count = 92317;
	#10 counter$count = 92318;
	#10 counter$count = 92319;
	#10 counter$count = 92320;
	#10 counter$count = 92321;
	#10 counter$count = 92322;
	#10 counter$count = 92323;
	#10 counter$count = 92324;
	#10 counter$count = 92325;
	#10 counter$count = 92326;
	#10 counter$count = 92327;
	#10 counter$count = 92328;
	#10 counter$count = 92329;
	#10 counter$count = 92330;
	#10 counter$count = 92331;
	#10 counter$count = 92332;
	#10 counter$count = 92333;
	#10 counter$count = 92334;
	#10 counter$count = 92335;
	#10 counter$count = 92336;
	#10 counter$count = 92337;
	#10 counter$count = 92338;
	#10 counter$count = 92339;
	#10 counter$count = 92340;
	#10 counter$count = 92341;
	#10 counter$count = 92342;
	#10 counter$count = 92343;
	#10 counter$count = 92344;
	#10 counter$count = 92345;
	#10 counter$count = 92346;
	#10 counter$count = 92347;
	#10 counter$count = 92348;
	#10 counter$count = 92349;
	#10 counter$count = 92350;
	#10 counter$count = 92351;
	#10 counter$count = 92352;
	#10 counter$count = 92353;
	#10 counter$count = 92354;
	#10 counter$count = 92355;
	#10 counter$count = 92356;
	#10 counter$count = 92357;
	#10 counter$count = 92358;
	#10 counter$count = 92359;
	#10 counter$count = 92360;
	#10 counter$count = 92361;
	#10 counter$count = 92362;
	#10 counter$count = 92363;
	#10 counter$count = 92364;
	#10 counter$count = 92365;
	#10 counter$count = 92366;
	#10 counter$count = 92367;
	#10 counter$count = 92368;
	#10 counter$count = 92369;
	#10 counter$count = 92370;
	#10 counter$count = 92371;
	#10 counter$count = 92372;
	#10 counter$count = 92373;
	#10 counter$count = 92374;
	#10 counter$count = 92375;
	#10 counter$count = 92376;
	#10 counter$count = 92377;
	#10 counter$count = 92378;
	#10 counter$count = 92379;
	#10 counter$count = 92380;
	#10 counter$count = 92381;
	#10 counter$count = 92382;
	#10 counter$count = 92383;
	#10 counter$count = 92384;
	#10 counter$count = 92385;
	#10 counter$count = 92386;
	#10 counter$count = 92387;
	#10 counter$count = 92388;
	#10 counter$count = 92389;
	#10 counter$count = 92390;
	#10 counter$count = 92391;
	#10 counter$count = 92392;
	#10 counter$count = 92393;
	#10 counter$count = 92394;
	#10 counter$count = 92395;
	#10 counter$count = 92396;
	#10 counter$count = 92397;
	#10 counter$count = 92398;
	#10 counter$count = 92399;
	#10 counter$count = 92400;
	#10 counter$count = 92401;
	#10 counter$count = 92402;
	#10 counter$count = 92403;
	#10 counter$count = 92404;
	#10 counter$count = 92405;
	#10 counter$count = 92406;
	#10 counter$count = 92407;
	#10 counter$count = 92408;
	#10 counter$count = 92409;
	#10 counter$count = 92410;
	#10 counter$count = 92411;
	#10 counter$count = 92412;
	#10 counter$count = 92413;
	#10 counter$count = 92414;
	#10 counter$count = 92415;
	#10 counter$count = 92416;
	#10 counter$count = 92417;
	#10 counter$count = 92418;
	#10 counter$count = 92419;
	#10 counter$count = 92420;
	#10 counter$count = 92421;
	#10 counter$count = 92422;
	#10 counter$count = 92423;
	#10 counter$count = 92424;
	#10 counter$count = 92425;
	#10 counter$count = 92426;
	#10 counter$count = 92427;
	#10 counter$count = 92428;
	#10 counter$count = 92429;
	#10 counter$count = 92430;
	#10 counter$count = 92431;
	#10 counter$count = 92432;
	#10 counter$count = 92433;
	#10 counter$count = 92434;
	#10 counter$count = 92435;
	#10 counter$count = 92436;
	#10 counter$count = 92437;
	#10 counter$count = 92438;
	#10 counter$count = 92439;
	#10 counter$count = 92440;
	#10 counter$count = 92441;
	#10 counter$count = 92442;
	#10 counter$count = 92443;
	#10 counter$count = 92444;
	#10 counter$count = 92445;
	#10 counter$count = 92446;
	#10 counter$count = 92447;
	#10 counter$count = 92448;
	#10 counter$count = 92449;
	#10 counter$count = 92450;
	#10 counter$count = 92451;
	#10 counter$count = 92452;
	#10 counter$count = 92453;
	#10 counter$count = 92454;
	#10 counter$count = 92455;
	#10 counter$count = 92456;
	#10 counter$count = 92457;
	#10 counter$count = 92458;
	#10 counter$count = 92459;
	#10 counter$count = 92460;
	#10 counter$count = 92461;
	#10 counter$count = 92462;
	#10 counter$count = 92463;
	#10 counter$count = 92464;
	#10 counter$count = 92465;
	#10 counter$count = 92466;
	#10 counter$count = 92467;
	#10 counter$count = 92468;
	#10 counter$count = 92469;
	#10 counter$count = 92470;
	#10 counter$count = 92471;
	#10 counter$count = 92472;
	#10 counter$count = 92473;
	#10 counter$count = 92474;
	#10 counter$count = 92475;
	#10 counter$count = 92476;
	#10 counter$count = 92477;
	#10 counter$count = 92478;
	#10 counter$count = 92479;
	#10 counter$count = 92480;
	#10 counter$count = 92481;
	#10 counter$count = 92482;
	#10 counter$count = 92483;
	#10 counter$count = 92484;
	#10 counter$count = 92485;
	#10 counter$count = 92486;
	#10 counter$count = 92487;
	#10 counter$count = 92488;
	#10 counter$count = 92489;
	#10 counter$count = 92490;
	#10 counter$count = 92491;
	#10 counter$count = 92492;
	#10 counter$count = 92493;
	#10 counter$count = 92494;
	#10 counter$count = 92495;
	#10 counter$count = 92496;
	#10 counter$count = 92497;
	#10 counter$count = 92498;
	#10 counter$count = 92499;
	#10 counter$count = 92500;
	#10 counter$count = 92501;
	#10 counter$count = 92502;
	#10 counter$count = 92503;
	#10 counter$count = 92504;
	#10 counter$count = 92505;
	#10 counter$count = 92506;
	#10 counter$count = 92507;
	#10 counter$count = 92508;
	#10 counter$count = 92509;
	#10 counter$count = 92510;
	#10 counter$count = 92511;
	#10 counter$count = 92512;
	#10 counter$count = 92513;
	#10 counter$count = 92514;
	#10 counter$count = 92515;
	#10 counter$count = 92516;
	#10 counter$count = 92517;
	#10 counter$count = 92518;
	#10 counter$count = 92519;
	#10 counter$count = 92520;
	#10 counter$count = 92521;
	#10 counter$count = 92522;
	#10 counter$count = 92523;
	#10 counter$count = 92524;
	#10 counter$count = 92525;
	#10 counter$count = 92526;
	#10 counter$count = 92527;
	#10 counter$count = 92528;
	#10 counter$count = 92529;
	#10 counter$count = 92530;
	#10 counter$count = 92531;
	#10 counter$count = 92532;
	#10 counter$count = 92533;
	#10 counter$count = 92534;
	#10 counter$count = 92535;
	#10 counter$count = 92536;
	#10 counter$count = 92537;
	#10 counter$count = 92538;
	#10 counter$count = 92539;
	#10 counter$count = 92540;
	#10 counter$count = 92541;
	#10 counter$count = 92542;
	#10 counter$count = 92543;
	#10 counter$count = 92544;
	#10 counter$count = 92545;
	#10 counter$count = 92546;
	#10 counter$count = 92547;
	#10 counter$count = 92548;
	#10 counter$count = 92549;
	#10 counter$count = 92550;
	#10 counter$count = 92551;
	#10 counter$count = 92552;
	#10 counter$count = 92553;
	#10 counter$count = 92554;
	#10 counter$count = 92555;
	#10 counter$count = 92556;
	#10 counter$count = 92557;
	#10 counter$count = 92558;
	#10 counter$count = 92559;
	#10 counter$count = 92560;
	#10 counter$count = 92561;
	#10 counter$count = 92562;
	#10 counter$count = 92563;
	#10 counter$count = 92564;
	#10 counter$count = 92565;
	#10 counter$count = 92566;
	#10 counter$count = 92567;
	#10 counter$count = 92568;
	#10 counter$count = 92569;
	#10 counter$count = 92570;
	#10 counter$count = 92571;
	#10 counter$count = 92572;
	#10 counter$count = 92573;
	#10 counter$count = 92574;
	#10 counter$count = 92575;
	#10 counter$count = 92576;
	#10 counter$count = 92577;
	#10 counter$count = 92578;
	#10 counter$count = 92579;
	#10 counter$count = 92580;
	#10 counter$count = 92581;
	#10 counter$count = 92582;
	#10 counter$count = 92583;
	#10 counter$count = 92584;
	#10 counter$count = 92585;
	#10 counter$count = 92586;
	#10 counter$count = 92587;
	#10 counter$count = 92588;
	#10 counter$count = 92589;
	#10 counter$count = 92590;
	#10 counter$count = 92591;
	#10 counter$count = 92592;
	#10 counter$count = 92593;
	#10 counter$count = 92594;
	#10 counter$count = 92595;
	#10 counter$count = 92596;
	#10 counter$count = 92597;
	#10 counter$count = 92598;
	#10 counter$count = 92599;
	#10 counter$count = 92600;
	#10 counter$count = 92601;
	#10 counter$count = 92602;
	#10 counter$count = 92603;
	#10 counter$count = 92604;
	#10 counter$count = 92605;
	#10 counter$count = 92606;
	#10 counter$count = 92607;
	#10 counter$count = 92608;
	#10 counter$count = 92609;
	#10 counter$count = 92610;
	#10 counter$count = 92611;
	#10 counter$count = 92612;
	#10 counter$count = 92613;
	#10 counter$count = 92614;
	#10 counter$count = 92615;
	#10 counter$count = 92616;
	#10 counter$count = 92617;
	#10 counter$count = 92618;
	#10 counter$count = 92619;
	#10 counter$count = 92620;
	#10 counter$count = 92621;
	#10 counter$count = 92622;
	#10 counter$count = 92623;
	#10 counter$count = 92624;
	#10 counter$count = 92625;
	#10 counter$count = 92626;
	#10 counter$count = 92627;
	#10 counter$count = 92628;
	#10 counter$count = 92629;
	#10 counter$count = 92630;
	#10 counter$count = 92631;
	#10 counter$count = 92632;
	#10 counter$count = 92633;
	#10 counter$count = 92634;
	#10 counter$count = 92635;
	#10 counter$count = 92636;
	#10 counter$count = 92637;
	#10 counter$count = 92638;
	#10 counter$count = 92639;
	#10 counter$count = 92640;
	#10 counter$count = 92641;
	#10 counter$count = 92642;
	#10 counter$count = 92643;
	#10 counter$count = 92644;
	#10 counter$count = 92645;
	#10 counter$count = 92646;
	#10 counter$count = 92647;
	#10 counter$count = 92648;
	#10 counter$count = 92649;
	#10 counter$count = 92650;
	#10 counter$count = 92651;
	#10 counter$count = 92652;
	#10 counter$count = 92653;
	#10 counter$count = 92654;
	#10 counter$count = 92655;
	#10 counter$count = 92656;
	#10 counter$count = 92657;
	#10 counter$count = 92658;
	#10 counter$count = 92659;
	#10 counter$count = 92660;
	#10 counter$count = 92661;
	#10 counter$count = 92662;
	#10 counter$count = 92663;
	#10 counter$count = 92664;
	#10 counter$count = 92665;
	#10 counter$count = 92666;
	#10 counter$count = 92667;
	#10 counter$count = 92668;
	#10 counter$count = 92669;
	#10 counter$count = 92670;
	#10 counter$count = 92671;
	#10 counter$count = 92672;
	#10 counter$count = 92673;
	#10 counter$count = 92674;
	#10 counter$count = 92675;
	#10 counter$count = 92676;
	#10 counter$count = 92677;
	#10 counter$count = 92678;
	#10 counter$count = 92679;
	#10 counter$count = 92680;
	#10 counter$count = 92681;
	#10 counter$count = 92682;
	#10 counter$count = 92683;
	#10 counter$count = 92684;
	#10 counter$count = 92685;
	#10 counter$count = 92686;
	#10 counter$count = 92687;
	#10 counter$count = 92688;
	#10 counter$count = 92689;
	#10 counter$count = 92690;
	#10 counter$count = 92691;
	#10 counter$count = 92692;
	#10 counter$count = 92693;
	#10 counter$count = 92694;
	#10 counter$count = 92695;
	#10 counter$count = 92696;
	#10 counter$count = 92697;
	#10 counter$count = 92698;
	#10 counter$count = 92699;
	#10 counter$count = 92700;
	#10 counter$count = 92701;
	#10 counter$count = 92702;
	#10 counter$count = 92703;
	#10 counter$count = 92704;
	#10 counter$count = 92705;
	#10 counter$count = 92706;
	#10 counter$count = 92707;
	#10 counter$count = 92708;
	#10 counter$count = 92709;
	#10 counter$count = 92710;
	#10 counter$count = 92711;
	#10 counter$count = 92712;
	#10 counter$count = 92713;
	#10 counter$count = 92714;
	#10 counter$count = 92715;
	#10 counter$count = 92716;
	#10 counter$count = 92717;
	#10 counter$count = 92718;
	#10 counter$count = 92719;
	#10 counter$count = 92720;
	#10 counter$count = 92721;
	#10 counter$count = 92722;
	#10 counter$count = 92723;
	#10 counter$count = 92724;
	#10 counter$count = 92725;
	#10 counter$count = 92726;
	#10 counter$count = 92727;
	#10 counter$count = 92728;
	#10 counter$count = 92729;
	#10 counter$count = 92730;
	#10 counter$count = 92731;
	#10 counter$count = 92732;
	#10 counter$count = 92733;
	#10 counter$count = 92734;
	#10 counter$count = 92735;
	#10 counter$count = 92736;
	#10 counter$count = 92737;
	#10 counter$count = 92738;
	#10 counter$count = 92739;
	#10 counter$count = 92740;
	#10 counter$count = 92741;
	#10 counter$count = 92742;
	#10 counter$count = 92743;
	#10 counter$count = 92744;
	#10 counter$count = 92745;
	#10 counter$count = 92746;
	#10 counter$count = 92747;
	#10 counter$count = 92748;
	#10 counter$count = 92749;
	#10 counter$count = 92750;
	#10 counter$count = 92751;
	#10 counter$count = 92752;
	#10 counter$count = 92753;
	#10 counter$count = 92754;
	#10 counter$count = 92755;
	#10 counter$count = 92756;
	#10 counter$count = 92757;
	#10 counter$count = 92758;
	#10 counter$count = 92759;
	#10 counter$count = 92760;
	#10 counter$count = 92761;
	#10 counter$count = 92762;
	#10 counter$count = 92763;
	#10 counter$count = 92764;
	#10 counter$count = 92765;
	#10 counter$count = 92766;
	#10 counter$count = 92767;
	#10 counter$count = 92768;
	#10 counter$count = 92769;
	#10 counter$count = 92770;
	#10 counter$count = 92771;
	#10 counter$count = 92772;
	#10 counter$count = 92773;
	#10 counter$count = 92774;
	#10 counter$count = 92775;
	#10 counter$count = 92776;
	#10 counter$count = 92777;
	#10 counter$count = 92778;
	#10 counter$count = 92779;
	#10 counter$count = 92780;
	#10 counter$count = 92781;
	#10 counter$count = 92782;
	#10 counter$count = 92783;
	#10 counter$count = 92784;
	#10 counter$count = 92785;
	#10 counter$count = 92786;
	#10 counter$count = 92787;
	#10 counter$count = 92788;
	#10 counter$count = 92789;
	#10 counter$count = 92790;
	#10 counter$count = 92791;
	#10 counter$count = 92792;
	#10 counter$count = 92793;
	#10 counter$count = 92794;
	#10 counter$count = 92795;
	#10 counter$count = 92796;
	#10 counter$count = 92797;
	#10 counter$count = 92798;
	#10 counter$count = 92799;
	#10 counter$count = 92800;
	#10 counter$count = 92801;
	#10 counter$count = 92802;
	#10 counter$count = 92803;
	#10 counter$count = 92804;
	#10 counter$count = 92805;
	#10 counter$count = 92806;
	#10 counter$count = 92807;
	#10 counter$count = 92808;
	#10 counter$count = 92809;
	#10 counter$count = 92810;
	#10 counter$count = 92811;
	#10 counter$count = 92812;
	#10 counter$count = 92813;
	#10 counter$count = 92814;
	#10 counter$count = 92815;
	#10 counter$count = 92816;
	#10 counter$count = 92817;
	#10 counter$count = 92818;
	#10 counter$count = 92819;
	#10 counter$count = 92820;
	#10 counter$count = 92821;
	#10 counter$count = 92822;
	#10 counter$count = 92823;
	#10 counter$count = 92824;
	#10 counter$count = 92825;
	#10 counter$count = 92826;
	#10 counter$count = 92827;
	#10 counter$count = 92828;
	#10 counter$count = 92829;
	#10 counter$count = 92830;
	#10 counter$count = 92831;
	#10 counter$count = 92832;
	#10 counter$count = 92833;
	#10 counter$count = 92834;
	#10 counter$count = 92835;
	#10 counter$count = 92836;
	#10 counter$count = 92837;
	#10 counter$count = 92838;
	#10 counter$count = 92839;
	#10 counter$count = 92840;
	#10 counter$count = 92841;
	#10 counter$count = 92842;
	#10 counter$count = 92843;
	#10 counter$count = 92844;
	#10 counter$count = 92845;
	#10 counter$count = 92846;
	#10 counter$count = 92847;
	#10 counter$count = 92848;
	#10 counter$count = 92849;
	#10 counter$count = 92850;
	#10 counter$count = 92851;
	#10 counter$count = 92852;
	#10 counter$count = 92853;
	#10 counter$count = 92854;
	#10 counter$count = 92855;
	#10 counter$count = 92856;
	#10 counter$count = 92857;
	#10 counter$count = 92858;
	#10 counter$count = 92859;
	#10 counter$count = 92860;
	#10 counter$count = 92861;
	#10 counter$count = 92862;
	#10 counter$count = 92863;
	#10 counter$count = 92864;
	#10 counter$count = 92865;
	#10 counter$count = 92866;
	#10 counter$count = 92867;
	#10 counter$count = 92868;
	#10 counter$count = 92869;
	#10 counter$count = 92870;
	#10 counter$count = 92871;
	#10 counter$count = 92872;
	#10 counter$count = 92873;
	#10 counter$count = 92874;
	#10 counter$count = 92875;
	#10 counter$count = 92876;
	#10 counter$count = 92877;
	#10 counter$count = 92878;
	#10 counter$count = 92879;
	#10 counter$count = 92880;
	#10 counter$count = 92881;
	#10 counter$count = 92882;
	#10 counter$count = 92883;
	#10 counter$count = 92884;
	#10 counter$count = 92885;
	#10 counter$count = 92886;
	#10 counter$count = 92887;
	#10 counter$count = 92888;
	#10 counter$count = 92889;
	#10 counter$count = 92890;
	#10 counter$count = 92891;
	#10 counter$count = 92892;
	#10 counter$count = 92893;
	#10 counter$count = 92894;
	#10 counter$count = 92895;
	#10 counter$count = 92896;
	#10 counter$count = 92897;
	#10 counter$count = 92898;
	#10 counter$count = 92899;
	#10 counter$count = 92900;
	#10 counter$count = 92901;
	#10 counter$count = 92902;
	#10 counter$count = 92903;
	#10 counter$count = 92904;
	#10 counter$count = 92905;
	#10 counter$count = 92906;
	#10 counter$count = 92907;
	#10 counter$count = 92908;
	#10 counter$count = 92909;
	#10 counter$count = 92910;
	#10 counter$count = 92911;
	#10 counter$count = 92912;
	#10 counter$count = 92913;
	#10 counter$count = 92914;
	#10 counter$count = 92915;
	#10 counter$count = 92916;
	#10 counter$count = 92917;
	#10 counter$count = 92918;
	#10 counter$count = 92919;
	#10 counter$count = 92920;
	#10 counter$count = 92921;
	#10 counter$count = 92922;
	#10 counter$count = 92923;
	#10 counter$count = 92924;
	#10 counter$count = 92925;
	#10 counter$count = 92926;
	#10 counter$count = 92927;
	#10 counter$count = 92928;
	#10 counter$count = 92929;
	#10 counter$count = 92930;
	#10 counter$count = 92931;
	#10 counter$count = 92932;
	#10 counter$count = 92933;
	#10 counter$count = 92934;
	#10 counter$count = 92935;
	#10 counter$count = 92936;
	#10 counter$count = 92937;
	#10 counter$count = 92938;
	#10 counter$count = 92939;
	#10 counter$count = 92940;
	#10 counter$count = 92941;
	#10 counter$count = 92942;
	#10 counter$count = 92943;
	#10 counter$count = 92944;
	#10 counter$count = 92945;
	#10 counter$count = 92946;
	#10 counter$count = 92947;
	#10 counter$count = 92948;
	#10 counter$count = 92949;
	#10 counter$count = 92950;
	#10 counter$count = 92951;
	#10 counter$count = 92952;
	#10 counter$count = 92953;
	#10 counter$count = 92954;
	#10 counter$count = 92955;
	#10 counter$count = 92956;
	#10 counter$count = 92957;
	#10 counter$count = 92958;
	#10 counter$count = 92959;
	#10 counter$count = 92960;
	#10 counter$count = 92961;
	#10 counter$count = 92962;
	#10 counter$count = 92963;
	#10 counter$count = 92964;
	#10 counter$count = 92965;
	#10 counter$count = 92966;
	#10 counter$count = 92967;
	#10 counter$count = 92968;
	#10 counter$count = 92969;
	#10 counter$count = 92970;
	#10 counter$count = 92971;
	#10 counter$count = 92972;
	#10 counter$count = 92973;
	#10 counter$count = 92974;
	#10 counter$count = 92975;
	#10 counter$count = 92976;
	#10 counter$count = 92977;
	#10 counter$count = 92978;
	#10 counter$count = 92979;
	#10 counter$count = 92980;
	#10 counter$count = 92981;
	#10 counter$count = 92982;
	#10 counter$count = 92983;
	#10 counter$count = 92984;
	#10 counter$count = 92985;
	#10 counter$count = 92986;
	#10 counter$count = 92987;
	#10 counter$count = 92988;
	#10 counter$count = 92989;
	#10 counter$count = 92990;
	#10 counter$count = 92991;
	#10 counter$count = 92992;
	#10 counter$count = 92993;
	#10 counter$count = 92994;
	#10 counter$count = 92995;
	#10 counter$count = 92996;
	#10 counter$count = 92997;
	#10 counter$count = 92998;
	#10 counter$count = 92999;
	#10 counter$count = 93000;
	#10 counter$count = 93001;
	#10 counter$count = 93002;
	#10 counter$count = 93003;
	#10 counter$count = 93004;
	#10 counter$count = 93005;
	#10 counter$count = 93006;
	#10 counter$count = 93007;
	#10 counter$count = 93008;
	#10 counter$count = 93009;
	#10 counter$count = 93010;
	#10 counter$count = 93011;
	#10 counter$count = 93012;
	#10 counter$count = 93013;
	#10 counter$count = 93014;
	#10 counter$count = 93015;
	#10 counter$count = 93016;
	#10 counter$count = 93017;
	#10 counter$count = 93018;
	#10 counter$count = 93019;
	#10 counter$count = 93020;
	#10 counter$count = 93021;
	#10 counter$count = 93022;
	#10 counter$count = 93023;
	#10 counter$count = 93024;
	#10 counter$count = 93025;
	#10 counter$count = 93026;
	#10 counter$count = 93027;
	#10 counter$count = 93028;
	#10 counter$count = 93029;
	#10 counter$count = 93030;
	#10 counter$count = 93031;
	#10 counter$count = 93032;
	#10 counter$count = 93033;
	#10 counter$count = 93034;
	#10 counter$count = 93035;
	#10 counter$count = 93036;
	#10 counter$count = 93037;
	#10 counter$count = 93038;
	#10 counter$count = 93039;
	#10 counter$count = 93040;
	#10 counter$count = 93041;
	#10 counter$count = 93042;
	#10 counter$count = 93043;
	#10 counter$count = 93044;
	#10 counter$count = 93045;
	#10 counter$count = 93046;
	#10 counter$count = 93047;
	#10 counter$count = 93048;
	#10 counter$count = 93049;
	#10 counter$count = 93050;
	#10 counter$count = 93051;
	#10 counter$count = 93052;
	#10 counter$count = 93053;
	#10 counter$count = 93054;
	#10 counter$count = 93055;
	#10 counter$count = 93056;
	#10 counter$count = 93057;
	#10 counter$count = 93058;
	#10 counter$count = 93059;
	#10 counter$count = 93060;
	#10 counter$count = 93061;
	#10 counter$count = 93062;
	#10 counter$count = 93063;
	#10 counter$count = 93064;
	#10 counter$count = 93065;
	#10 counter$count = 93066;
	#10 counter$count = 93067;
	#10 counter$count = 93068;
	#10 counter$count = 93069;
	#10 counter$count = 93070;
	#10 counter$count = 93071;
	#10 counter$count = 93072;
	#10 counter$count = 93073;
	#10 counter$count = 93074;
	#10 counter$count = 93075;
	#10 counter$count = 93076;
	#10 counter$count = 93077;
	#10 counter$count = 93078;
	#10 counter$count = 93079;
	#10 counter$count = 93080;
	#10 counter$count = 93081;
	#10 counter$count = 93082;
	#10 counter$count = 93083;
	#10 counter$count = 93084;
	#10 counter$count = 93085;
	#10 counter$count = 93086;
	#10 counter$count = 93087;
	#10 counter$count = 93088;
	#10 counter$count = 93089;
	#10 counter$count = 93090;
	#10 counter$count = 93091;
	#10 counter$count = 93092;
	#10 counter$count = 93093;
	#10 counter$count = 93094;
	#10 counter$count = 93095;
	#10 counter$count = 93096;
	#10 counter$count = 93097;
	#10 counter$count = 93098;
	#10 counter$count = 93099;
	#10 counter$count = 93100;
	#10 counter$count = 93101;
	#10 counter$count = 93102;
	#10 counter$count = 93103;
	#10 counter$count = 93104;
	#10 counter$count = 93105;
	#10 counter$count = 93106;
	#10 counter$count = 93107;
	#10 counter$count = 93108;
	#10 counter$count = 93109;
	#10 counter$count = 93110;
	#10 counter$count = 93111;
	#10 counter$count = 93112;
	#10 counter$count = 93113;
	#10 counter$count = 93114;
	#10 counter$count = 93115;
	#10 counter$count = 93116;
	#10 counter$count = 93117;
	#10 counter$count = 93118;
	#10 counter$count = 93119;
	#10 counter$count = 93120;
	#10 counter$count = 93121;
	#10 counter$count = 93122;
	#10 counter$count = 93123;
	#10 counter$count = 93124;
	#10 counter$count = 93125;
	#10 counter$count = 93126;
	#10 counter$count = 93127;
	#10 counter$count = 93128;
	#10 counter$count = 93129;
	#10 counter$count = 93130;
	#10 counter$count = 93131;
	#10 counter$count = 93132;
	#10 counter$count = 93133;
	#10 counter$count = 93134;
	#10 counter$count = 93135;
	#10 counter$count = 93136;
	#10 counter$count = 93137;
	#10 counter$count = 93138;
	#10 counter$count = 93139;
	#10 counter$count = 93140;
	#10 counter$count = 93141;
	#10 counter$count = 93142;
	#10 counter$count = 93143;
	#10 counter$count = 93144;
	#10 counter$count = 93145;
	#10 counter$count = 93146;
	#10 counter$count = 93147;
	#10 counter$count = 93148;
	#10 counter$count = 93149;
	#10 counter$count = 93150;
	#10 counter$count = 93151;
	#10 counter$count = 93152;
	#10 counter$count = 93153;
	#10 counter$count = 93154;
	#10 counter$count = 93155;
	#10 counter$count = 93156;
	#10 counter$count = 93157;
	#10 counter$count = 93158;
	#10 counter$count = 93159;
	#10 counter$count = 93160;
	#10 counter$count = 93161;
	#10 counter$count = 93162;
	#10 counter$count = 93163;
	#10 counter$count = 93164;
	#10 counter$count = 93165;
	#10 counter$count = 93166;
	#10 counter$count = 93167;
	#10 counter$count = 93168;
	#10 counter$count = 93169;
	#10 counter$count = 93170;
	#10 counter$count = 93171;
	#10 counter$count = 93172;
	#10 counter$count = 93173;
	#10 counter$count = 93174;
	#10 counter$count = 93175;
	#10 counter$count = 93176;
	#10 counter$count = 93177;
	#10 counter$count = 93178;
	#10 counter$count = 93179;
	#10 counter$count = 93180;
	#10 counter$count = 93181;
	#10 counter$count = 93182;
	#10 counter$count = 93183;
	#10 counter$count = 93184;
	#10 counter$count = 93185;
	#10 counter$count = 93186;
	#10 counter$count = 93187;
	#10 counter$count = 93188;
	#10 counter$count = 93189;
	#10 counter$count = 93190;
	#10 counter$count = 93191;
	#10 counter$count = 93192;
	#10 counter$count = 93193;
	#10 counter$count = 93194;
	#10 counter$count = 93195;
	#10 counter$count = 93196;
	#10 counter$count = 93197;
	#10 counter$count = 93198;
	#10 counter$count = 93199;
	#10 counter$count = 93200;
	#10 counter$count = 93201;
	#10 counter$count = 93202;
	#10 counter$count = 93203;
	#10 counter$count = 93204;
	#10 counter$count = 93205;
	#10 counter$count = 93206;
	#10 counter$count = 93207;
	#10 counter$count = 93208;
	#10 counter$count = 93209;
	#10 counter$count = 93210;
	#10 counter$count = 93211;
	#10 counter$count = 93212;
	#10 counter$count = 93213;
	#10 counter$count = 93214;
	#10 counter$count = 93215;
	#10 counter$count = 93216;
	#10 counter$count = 93217;
	#10 counter$count = 93218;
	#10 counter$count = 93219;
	#10 counter$count = 93220;
	#10 counter$count = 93221;
	#10 counter$count = 93222;
	#10 counter$count = 93223;
	#10 counter$count = 93224;
	#10 counter$count = 93225;
	#10 counter$count = 93226;
	#10 counter$count = 93227;
	#10 counter$count = 93228;
	#10 counter$count = 93229;
	#10 counter$count = 93230;
	#10 counter$count = 93231;
	#10 counter$count = 93232;
	#10 counter$count = 93233;
	#10 counter$count = 93234;
	#10 counter$count = 93235;
	#10 counter$count = 93236;
	#10 counter$count = 93237;
	#10 counter$count = 93238;
	#10 counter$count = 93239;
	#10 counter$count = 93240;
	#10 counter$count = 93241;
	#10 counter$count = 93242;
	#10 counter$count = 93243;
	#10 counter$count = 93244;
	#10 counter$count = 93245;
	#10 counter$count = 93246;
	#10 counter$count = 93247;
	#10 counter$count = 93248;
	#10 counter$count = 93249;
	#10 counter$count = 93250;
	#10 counter$count = 93251;
	#10 counter$count = 93252;
	#10 counter$count = 93253;
	#10 counter$count = 93254;
	#10 counter$count = 93255;
	#10 counter$count = 93256;
	#10 counter$count = 93257;
	#10 counter$count = 93258;
	#10 counter$count = 93259;
	#10 counter$count = 93260;
	#10 counter$count = 93261;
	#10 counter$count = 93262;
	#10 counter$count = 93263;
	#10 counter$count = 93264;
	#10 counter$count = 93265;
	#10 counter$count = 93266;
	#10 counter$count = 93267;
	#10 counter$count = 93268;
	#10 counter$count = 93269;
	#10 counter$count = 93270;
	#10 counter$count = 93271;
	#10 counter$count = 93272;
	#10 counter$count = 93273;
	#10 counter$count = 93274;
	#10 counter$count = 93275;
	#10 counter$count = 93276;
	#10 counter$count = 93277;
	#10 counter$count = 93278;
	#10 counter$count = 93279;
	#10 counter$count = 93280;
	#10 counter$count = 93281;
	#10 counter$count = 93282;
	#10 counter$count = 93283;
	#10 counter$count = 93284;
	#10 counter$count = 93285;
	#10 counter$count = 93286;
	#10 counter$count = 93287;
	#10 counter$count = 93288;
	#10 counter$count = 93289;
	#10 counter$count = 93290;
	#10 counter$count = 93291;
	#10 counter$count = 93292;
	#10 counter$count = 93293;
	#10 counter$count = 93294;
	#10 counter$count = 93295;
	#10 counter$count = 93296;
	#10 counter$count = 93297;
	#10 counter$count = 93298;
	#10 counter$count = 93299;
	#10 counter$count = 93300;
	#10 counter$count = 93301;
	#10 counter$count = 93302;
	#10 counter$count = 93303;
	#10 counter$count = 93304;
	#10 counter$count = 93305;
	#10 counter$count = 93306;
	#10 counter$count = 93307;
	#10 counter$count = 93308;
	#10 counter$count = 93309;
	#10 counter$count = 93310;
	#10 counter$count = 93311;
	#10 counter$count = 93312;
	#10 counter$count = 93313;
	#10 counter$count = 93314;
	#10 counter$count = 93315;
	#10 counter$count = 93316;
	#10 counter$count = 93317;
	#10 counter$count = 93318;
	#10 counter$count = 93319;
	#10 counter$count = 93320;
	#10 counter$count = 93321;
	#10 counter$count = 93322;
	#10 counter$count = 93323;
	#10 counter$count = 93324;
	#10 counter$count = 93325;
	#10 counter$count = 93326;
	#10 counter$count = 93327;
	#10 counter$count = 93328;
	#10 counter$count = 93329;
	#10 counter$count = 93330;
	#10 counter$count = 93331;
	#10 counter$count = 93332;
	#10 counter$count = 93333;
	#10 counter$count = 93334;
	#10 counter$count = 93335;
	#10 counter$count = 93336;
	#10 counter$count = 93337;
	#10 counter$count = 93338;
	#10 counter$count = 93339;
	#10 counter$count = 93340;
	#10 counter$count = 93341;
	#10 counter$count = 93342;
	#10 counter$count = 93343;
	#10 counter$count = 93344;
	#10 counter$count = 93345;
	#10 counter$count = 93346;
	#10 counter$count = 93347;
	#10 counter$count = 93348;
	#10 counter$count = 93349;
	#10 counter$count = 93350;
	#10 counter$count = 93351;
	#10 counter$count = 93352;
	#10 counter$count = 93353;
	#10 counter$count = 93354;
	#10 counter$count = 93355;
	#10 counter$count = 93356;
	#10 counter$count = 93357;
	#10 counter$count = 93358;
	#10 counter$count = 93359;
	#10 counter$count = 93360;
	#10 counter$count = 93361;
	#10 counter$count = 93362;
	#10 counter$count = 93363;
	#10 counter$count = 93364;
	#10 counter$count = 93365;
	#10 counter$count = 93366;
	#10 counter$count = 93367;
	#10 counter$count = 93368;
	#10 counter$count = 93369;
	#10 counter$count = 93370;
	#10 counter$count = 93371;
	#10 counter$count = 93372;
	#10 counter$count = 93373;
	#10 counter$count = 93374;
	#10 counter$count = 93375;
	#10 counter$count = 93376;
	#10 counter$count = 93377;
	#10 counter$count = 93378;
	#10 counter$count = 93379;
	#10 counter$count = 93380;
	#10 counter$count = 93381;
	#10 counter$count = 93382;
	#10 counter$count = 93383;
	#10 counter$count = 93384;
	#10 counter$count = 93385;
	#10 counter$count = 93386;
	#10 counter$count = 93387;
	#10 counter$count = 93388;
	#10 counter$count = 93389;
	#10 counter$count = 93390;
	#10 counter$count = 93391;
	#10 counter$count = 93392;
	#10 counter$count = 93393;
	#10 counter$count = 93394;
	#10 counter$count = 93395;
	#10 counter$count = 93396;
	#10 counter$count = 93397;
	#10 counter$count = 93398;
	#10 counter$count = 93399;
	#10 counter$count = 93400;
	#10 counter$count = 93401;
	#10 counter$count = 93402;
	#10 counter$count = 93403;
	#10 counter$count = 93404;
	#10 counter$count = 93405;
	#10 counter$count = 93406;
	#10 counter$count = 93407;
	#10 counter$count = 93408;
	#10 counter$count = 93409;
	#10 counter$count = 93410;
	#10 counter$count = 93411;
	#10 counter$count = 93412;
	#10 counter$count = 93413;
	#10 counter$count = 93414;
	#10 counter$count = 93415;
	#10 counter$count = 93416;
	#10 counter$count = 93417;
	#10 counter$count = 93418;
	#10 counter$count = 93419;
	#10 counter$count = 93420;
	#10 counter$count = 93421;
	#10 counter$count = 93422;
	#10 counter$count = 93423;
	#10 counter$count = 93424;
	#10 counter$count = 93425;
	#10 counter$count = 93426;
	#10 counter$count = 93427;
	#10 counter$count = 93428;
	#10 counter$count = 93429;
	#10 counter$count = 93430;
	#10 counter$count = 93431;
	#10 counter$count = 93432;
	#10 counter$count = 93433;
	#10 counter$count = 93434;
	#10 counter$count = 93435;
	#10 counter$count = 93436;
	#10 counter$count = 93437;
	#10 counter$count = 93438;
	#10 counter$count = 93439;
	#10 counter$count = 93440;
	#10 counter$count = 93441;
	#10 counter$count = 93442;
	#10 counter$count = 93443;
	#10 counter$count = 93444;
	#10 counter$count = 93445;
	#10 counter$count = 93446;
	#10 counter$count = 93447;
	#10 counter$count = 93448;
	#10 counter$count = 93449;
	#10 counter$count = 93450;
	#10 counter$count = 93451;
	#10 counter$count = 93452;
	#10 counter$count = 93453;
	#10 counter$count = 93454;
	#10 counter$count = 93455;
	#10 counter$count = 93456;
	#10 counter$count = 93457;
	#10 counter$count = 93458;
	#10 counter$count = 93459;
	#10 counter$count = 93460;
	#10 counter$count = 93461;
	#10 counter$count = 93462;
	#10 counter$count = 93463;
	#10 counter$count = 93464;
	#10 counter$count = 93465;
	#10 counter$count = 93466;
	#10 counter$count = 93467;
	#10 counter$count = 93468;
	#10 counter$count = 93469;
	#10 counter$count = 93470;
	#10 counter$count = 93471;
	#10 counter$count = 93472;
	#10 counter$count = 93473;
	#10 counter$count = 93474;
	#10 counter$count = 93475;
	#10 counter$count = 93476;
	#10 counter$count = 93477;
	#10 counter$count = 93478;
	#10 counter$count = 93479;
	#10 counter$count = 93480;
	#10 counter$count = 93481;
	#10 counter$count = 93482;
	#10 counter$count = 93483;
	#10 counter$count = 93484;
	#10 counter$count = 93485;
	#10 counter$count = 93486;
	#10 counter$count = 93487;
	#10 counter$count = 93488;
	#10 counter$count = 93489;
	#10 counter$count = 93490;
	#10 counter$count = 93491;
	#10 counter$count = 93492;
	#10 counter$count = 93493;
	#10 counter$count = 93494;
	#10 counter$count = 93495;
	#10 counter$count = 93496;
	#10 counter$count = 93497;
	#10 counter$count = 93498;
	#10 counter$count = 93499;
	#10 counter$count = 93500;
	#10 counter$count = 93501;
	#10 counter$count = 93502;
	#10 counter$count = 93503;
	#10 counter$count = 93504;
	#10 counter$count = 93505;
	#10 counter$count = 93506;
	#10 counter$count = 93507;
	#10 counter$count = 93508;
	#10 counter$count = 93509;
	#10 counter$count = 93510;
	#10 counter$count = 93511;
	#10 counter$count = 93512;
	#10 counter$count = 93513;
	#10 counter$count = 93514;
	#10 counter$count = 93515;
	#10 counter$count = 93516;
	#10 counter$count = 93517;
	#10 counter$count = 93518;
	#10 counter$count = 93519;
	#10 counter$count = 93520;
	#10 counter$count = 93521;
	#10 counter$count = 93522;
	#10 counter$count = 93523;
	#10 counter$count = 93524;
	#10 counter$count = 93525;
	#10 counter$count = 93526;
	#10 counter$count = 93527;
	#10 counter$count = 93528;
	#10 counter$count = 93529;
	#10 counter$count = 93530;
	#10 counter$count = 93531;
	#10 counter$count = 93532;
	#10 counter$count = 93533;
	#10 counter$count = 93534;
	#10 counter$count = 93535;
	#10 counter$count = 93536;
	#10 counter$count = 93537;
	#10 counter$count = 93538;
	#10 counter$count = 93539;
	#10 counter$count = 93540;
	#10 counter$count = 93541;
	#10 counter$count = 93542;
	#10 counter$count = 93543;
	#10 counter$count = 93544;
	#10 counter$count = 93545;
	#10 counter$count = 93546;
	#10 counter$count = 93547;
	#10 counter$count = 93548;
	#10 counter$count = 93549;
	#10 counter$count = 93550;
	#10 counter$count = 93551;
	#10 counter$count = 93552;
	#10 counter$count = 93553;
	#10 counter$count = 93554;
	#10 counter$count = 93555;
	#10 counter$count = 93556;
	#10 counter$count = 93557;
	#10 counter$count = 93558;
	#10 counter$count = 93559;
	#10 counter$count = 93560;
	#10 counter$count = 93561;
	#10 counter$count = 93562;
	#10 counter$count = 93563;
	#10 counter$count = 93564;
	#10 counter$count = 93565;
	#10 counter$count = 93566;
	#10 counter$count = 93567;
	#10 counter$count = 93568;
	#10 counter$count = 93569;
	#10 counter$count = 93570;
	#10 counter$count = 93571;
	#10 counter$count = 93572;
	#10 counter$count = 93573;
	#10 counter$count = 93574;
	#10 counter$count = 93575;
	#10 counter$count = 93576;
	#10 counter$count = 93577;
	#10 counter$count = 93578;
	#10 counter$count = 93579;
	#10 counter$count = 93580;
	#10 counter$count = 93581;
	#10 counter$count = 93582;
	#10 counter$count = 93583;
	#10 counter$count = 93584;
	#10 counter$count = 93585;
	#10 counter$count = 93586;
	#10 counter$count = 93587;
	#10 counter$count = 93588;
	#10 counter$count = 93589;
	#10 counter$count = 93590;
	#10 counter$count = 93591;
	#10 counter$count = 93592;
	#10 counter$count = 93593;
	#10 counter$count = 93594;
	#10 counter$count = 93595;
	#10 counter$count = 93596;
	#10 counter$count = 93597;
	#10 counter$count = 93598;
	#10 counter$count = 93599;
	#10 counter$count = 93600;
	#10 counter$count = 93601;
	#10 counter$count = 93602;
	#10 counter$count = 93603;
	#10 counter$count = 93604;
	#10 counter$count = 93605;
	#10 counter$count = 93606;
	#10 counter$count = 93607;
	#10 counter$count = 93608;
	#10 counter$count = 93609;
	#10 counter$count = 93610;
	#10 counter$count = 93611;
	#10 counter$count = 93612;
	#10 counter$count = 93613;
	#10 counter$count = 93614;
	#10 counter$count = 93615;
	#10 counter$count = 93616;
	#10 counter$count = 93617;
	#10 counter$count = 93618;
	#10 counter$count = 93619;
	#10 counter$count = 93620;
	#10 counter$count = 93621;
	#10 counter$count = 93622;
	#10 counter$count = 93623;
	#10 counter$count = 93624;
	#10 counter$count = 93625;
	#10 counter$count = 93626;
	#10 counter$count = 93627;
	#10 counter$count = 93628;
	#10 counter$count = 93629;
	#10 counter$count = 93630;
	#10 counter$count = 93631;
	#10 counter$count = 93632;
	#10 counter$count = 93633;
	#10 counter$count = 93634;
	#10 counter$count = 93635;
	#10 counter$count = 93636;
	#10 counter$count = 93637;
	#10 counter$count = 93638;
	#10 counter$count = 93639;
	#10 counter$count = 93640;
	#10 counter$count = 93641;
	#10 counter$count = 93642;
	#10 counter$count = 93643;
	#10 counter$count = 93644;
	#10 counter$count = 93645;
	#10 counter$count = 93646;
	#10 counter$count = 93647;
	#10 counter$count = 93648;
	#10 counter$count = 93649;
	#10 counter$count = 93650;
	#10 counter$count = 93651;
	#10 counter$count = 93652;
	#10 counter$count = 93653;
	#10 counter$count = 93654;
	#10 counter$count = 93655;
	#10 counter$count = 93656;
	#10 counter$count = 93657;
	#10 counter$count = 93658;
	#10 counter$count = 93659;
	#10 counter$count = 93660;
	#10 counter$count = 93661;
	#10 counter$count = 93662;
	#10 counter$count = 93663;
	#10 counter$count = 93664;
	#10 counter$count = 93665;
	#10 counter$count = 93666;
	#10 counter$count = 93667;
	#10 counter$count = 93668;
	#10 counter$count = 93669;
	#10 counter$count = 93670;
	#10 counter$count = 93671;
	#10 counter$count = 93672;
	#10 counter$count = 93673;
	#10 counter$count = 93674;
	#10 counter$count = 93675;
	#10 counter$count = 93676;
	#10 counter$count = 93677;
	#10 counter$count = 93678;
	#10 counter$count = 93679;
	#10 counter$count = 93680;
	#10 counter$count = 93681;
	#10 counter$count = 93682;
	#10 counter$count = 93683;
	#10 counter$count = 93684;
	#10 counter$count = 93685;
	#10 counter$count = 93686;
	#10 counter$count = 93687;
	#10 counter$count = 93688;
	#10 counter$count = 93689;
	#10 counter$count = 93690;
	#10 counter$count = 93691;
	#10 counter$count = 93692;
	#10 counter$count = 93693;
	#10 counter$count = 93694;
	#10 counter$count = 93695;
	#10 counter$count = 93696;
	#10 counter$count = 93697;
	#10 counter$count = 93698;
	#10 counter$count = 93699;
	#10 counter$count = 93700;
	#10 counter$count = 93701;
	#10 counter$count = 93702;
	#10 counter$count = 93703;
	#10 counter$count = 93704;
	#10 counter$count = 93705;
	#10 counter$count = 93706;
	#10 counter$count = 93707;
	#10 counter$count = 93708;
	#10 counter$count = 93709;
	#10 counter$count = 93710;
	#10 counter$count = 93711;
	#10 counter$count = 93712;
	#10 counter$count = 93713;
	#10 counter$count = 93714;
	#10 counter$count = 93715;
	#10 counter$count = 93716;
	#10 counter$count = 93717;
	#10 counter$count = 93718;
	#10 counter$count = 93719;
	#10 counter$count = 93720;
	#10 counter$count = 93721;
	#10 counter$count = 93722;
	#10 counter$count = 93723;
	#10 counter$count = 93724;
	#10 counter$count = 93725;
	#10 counter$count = 93726;
	#10 counter$count = 93727;
	#10 counter$count = 93728;
	#10 counter$count = 93729;
	#10 counter$count = 93730;
	#10 counter$count = 93731;
	#10 counter$count = 93732;
	#10 counter$count = 93733;
	#10 counter$count = 93734;
	#10 counter$count = 93735;
	#10 counter$count = 93736;
	#10 counter$count = 93737;
	#10 counter$count = 93738;
	#10 counter$count = 93739;
	#10 counter$count = 93740;
	#10 counter$count = 93741;
	#10 counter$count = 93742;
	#10 counter$count = 93743;
	#10 counter$count = 93744;
	#10 counter$count = 93745;
	#10 counter$count = 93746;
	#10 counter$count = 93747;
	#10 counter$count = 93748;
	#10 counter$count = 93749;
	#10 counter$count = 93750;
	#10 counter$count = 93751;
	#10 counter$count = 93752;
	#10 counter$count = 93753;
	#10 counter$count = 93754;
	#10 counter$count = 93755;
	#10 counter$count = 93756;
	#10 counter$count = 93757;
	#10 counter$count = 93758;
	#10 counter$count = 93759;
	#10 counter$count = 93760;
	#10 counter$count = 93761;
	#10 counter$count = 93762;
	#10 counter$count = 93763;
	#10 counter$count = 93764;
	#10 counter$count = 93765;
	#10 counter$count = 93766;
	#10 counter$count = 93767;
	#10 counter$count = 93768;
	#10 counter$count = 93769;
	#10 counter$count = 93770;
	#10 counter$count = 93771;
	#10 counter$count = 93772;
	#10 counter$count = 93773;
	#10 counter$count = 93774;
	#10 counter$count = 93775;
	#10 counter$count = 93776;
	#10 counter$count = 93777;
	#10 counter$count = 93778;
	#10 counter$count = 93779;
	#10 counter$count = 93780;
	#10 counter$count = 93781;
	#10 counter$count = 93782;
	#10 counter$count = 93783;
	#10 counter$count = 93784;
	#10 counter$count = 93785;
	#10 counter$count = 93786;
	#10 counter$count = 93787;
	#10 counter$count = 93788;
	#10 counter$count = 93789;
	#10 counter$count = 93790;
	#10 counter$count = 93791;
	#10 counter$count = 93792;
	#10 counter$count = 93793;
	#10 counter$count = 93794;
	#10 counter$count = 93795;
	#10 counter$count = 93796;
	#10 counter$count = 93797;
	#10 counter$count = 93798;
	#10 counter$count = 93799;
	#10 counter$count = 93800;
	#10 counter$count = 93801;
	#10 counter$count = 93802;
	#10 counter$count = 93803;
	#10 counter$count = 93804;
	#10 counter$count = 93805;
	#10 counter$count = 93806;
	#10 counter$count = 93807;
	#10 counter$count = 93808;
	#10 counter$count = 93809;
	#10 counter$count = 93810;
	#10 counter$count = 93811;
	#10 counter$count = 93812;
	#10 counter$count = 93813;
	#10 counter$count = 93814;
	#10 counter$count = 93815;
	#10 counter$count = 93816;
	#10 counter$count = 93817;
	#10 counter$count = 93818;
	#10 counter$count = 93819;
	#10 counter$count = 93820;
	#10 counter$count = 93821;
	#10 counter$count = 93822;
	#10 counter$count = 93823;
	#10 counter$count = 93824;
	#10 counter$count = 93825;
	#10 counter$count = 93826;
	#10 counter$count = 93827;
	#10 counter$count = 93828;
	#10 counter$count = 93829;
	#10 counter$count = 93830;
	#10 counter$count = 93831;
	#10 counter$count = 93832;
	#10 counter$count = 93833;
	#10 counter$count = 93834;
	#10 counter$count = 93835;
	#10 counter$count = 93836;
	#10 counter$count = 93837;
	#10 counter$count = 93838;
	#10 counter$count = 93839;
	#10 counter$count = 93840;
	#10 counter$count = 93841;
	#10 counter$count = 93842;
	#10 counter$count = 93843;
	#10 counter$count = 93844;
	#10 counter$count = 93845;
	#10 counter$count = 93846;
	#10 counter$count = 93847;
	#10 counter$count = 93848;
	#10 counter$count = 93849;
	#10 counter$count = 93850;
	#10 counter$count = 93851;
	#10 counter$count = 93852;
	#10 counter$count = 93853;
	#10 counter$count = 93854;
	#10 counter$count = 93855;
	#10 counter$count = 93856;
	#10 counter$count = 93857;
	#10 counter$count = 93858;
	#10 counter$count = 93859;
	#10 counter$count = 93860;
	#10 counter$count = 93861;
	#10 counter$count = 93862;
	#10 counter$count = 93863;
	#10 counter$count = 93864;
	#10 counter$count = 93865;
	#10 counter$count = 93866;
	#10 counter$count = 93867;
	#10 counter$count = 93868;
	#10 counter$count = 93869;
	#10 counter$count = 93870;
	#10 counter$count = 93871;
	#10 counter$count = 93872;
	#10 counter$count = 93873;
	#10 counter$count = 93874;
	#10 counter$count = 93875;
	#10 counter$count = 93876;
	#10 counter$count = 93877;
	#10 counter$count = 93878;
	#10 counter$count = 93879;
	#10 counter$count = 93880;
	#10 counter$count = 93881;
	#10 counter$count = 93882;
	#10 counter$count = 93883;
	#10 counter$count = 93884;
	#10 counter$count = 93885;
	#10 counter$count = 93886;
	#10 counter$count = 93887;
	#10 counter$count = 93888;
	#10 counter$count = 93889;
	#10 counter$count = 93890;
	#10 counter$count = 93891;
	#10 counter$count = 93892;
	#10 counter$count = 93893;
	#10 counter$count = 93894;
	#10 counter$count = 93895;
	#10 counter$count = 93896;
	#10 counter$count = 93897;
	#10 counter$count = 93898;
	#10 counter$count = 93899;
	#10 counter$count = 93900;
	#10 counter$count = 93901;
	#10 counter$count = 93902;
	#10 counter$count = 93903;
	#10 counter$count = 93904;
	#10 counter$count = 93905;
	#10 counter$count = 93906;
	#10 counter$count = 93907;
	#10 counter$count = 93908;
	#10 counter$count = 93909;
	#10 counter$count = 93910;
	#10 counter$count = 93911;
	#10 counter$count = 93912;
	#10 counter$count = 93913;
	#10 counter$count = 93914;
	#10 counter$count = 93915;
	#10 counter$count = 93916;
	#10 counter$count = 93917;
	#10 counter$count = 93918;
	#10 counter$count = 93919;
	#10 counter$count = 93920;
	#10 counter$count = 93921;
	#10 counter$count = 93922;
	#10 counter$count = 93923;
	#10 counter$count = 93924;
	#10 counter$count = 93925;
	#10 counter$count = 93926;
	#10 counter$count = 93927;
	#10 counter$count = 93928;
	#10 counter$count = 93929;
	#10 counter$count = 93930;
	#10 counter$count = 93931;
	#10 counter$count = 93932;
	#10 counter$count = 93933;
	#10 counter$count = 93934;
	#10 counter$count = 93935;
	#10 counter$count = 93936;
	#10 counter$count = 93937;
	#10 counter$count = 93938;
	#10 counter$count = 93939;
	#10 counter$count = 93940;
	#10 counter$count = 93941;
	#10 counter$count = 93942;
	#10 counter$count = 93943;
	#10 counter$count = 93944;
	#10 counter$count = 93945;
	#10 counter$count = 93946;
	#10 counter$count = 93947;
	#10 counter$count = 93948;
	#10 counter$count = 93949;
	#10 counter$count = 93950;
	#10 counter$count = 93951;
	#10 counter$count = 93952;
	#10 counter$count = 93953;
	#10 counter$count = 93954;
	#10 counter$count = 93955;
	#10 counter$count = 93956;
	#10 counter$count = 93957;
	#10 counter$count = 93958;
	#10 counter$count = 93959;
	#10 counter$count = 93960;
	#10 counter$count = 93961;
	#10 counter$count = 93962;
	#10 counter$count = 93963;
	#10 counter$count = 93964;
	#10 counter$count = 93965;
	#10 counter$count = 93966;
	#10 counter$count = 93967;
	#10 counter$count = 93968;
	#10 counter$count = 93969;
	#10 counter$count = 93970;
	#10 counter$count = 93971;
	#10 counter$count = 93972;
	#10 counter$count = 93973;
	#10 counter$count = 93974;
	#10 counter$count = 93975;
	#10 counter$count = 93976;
	#10 counter$count = 93977;
	#10 counter$count = 93978;
	#10 counter$count = 93979;
	#10 counter$count = 93980;
	#10 counter$count = 93981;
	#10 counter$count = 93982;
	#10 counter$count = 93983;
	#10 counter$count = 93984;
	#10 counter$count = 93985;
	#10 counter$count = 93986;
	#10 counter$count = 93987;
	#10 counter$count = 93988;
	#10 counter$count = 93989;
	#10 counter$count = 93990;
	#10 counter$count = 93991;
	#10 counter$count = 93992;
	#10 counter$count = 93993;
	#10 counter$count = 93994;
	#10 counter$count = 93995;
	#10 counter$count = 93996;
	#10 counter$count = 93997;
	#10 counter$count = 93998;
	#10 counter$count = 93999;
	#10 counter$count = 94000;
	#10 counter$count = 94001;
	#10 counter$count = 94002;
	#10 counter$count = 94003;
	#10 counter$count = 94004;
	#10 counter$count = 94005;
	#10 counter$count = 94006;
	#10 counter$count = 94007;
	#10 counter$count = 94008;
	#10 counter$count = 94009;
	#10 counter$count = 94010;
	#10 counter$count = 94011;
	#10 counter$count = 94012;
	#10 counter$count = 94013;
	#10 counter$count = 94014;
	#10 counter$count = 94015;
	#10 counter$count = 94016;
	#10 counter$count = 94017;
	#10 counter$count = 94018;
	#10 counter$count = 94019;
	#10 counter$count = 94020;
	#10 counter$count = 94021;
	#10 counter$count = 94022;
	#10 counter$count = 94023;
	#10 counter$count = 94024;
	#10 counter$count = 94025;
	#10 counter$count = 94026;
	#10 counter$count = 94027;
	#10 counter$count = 94028;
	#10 counter$count = 94029;
	#10 counter$count = 94030;
	#10 counter$count = 94031;
	#10 counter$count = 94032;
	#10 counter$count = 94033;
	#10 counter$count = 94034;
	#10 counter$count = 94035;
	#10 counter$count = 94036;
	#10 counter$count = 94037;
	#10 counter$count = 94038;
	#10 counter$count = 94039;
	#10 counter$count = 94040;
	#10 counter$count = 94041;
	#10 counter$count = 94042;
	#10 counter$count = 94043;
	#10 counter$count = 94044;
	#10 counter$count = 94045;
	#10 counter$count = 94046;
	#10 counter$count = 94047;
	#10 counter$count = 94048;
	#10 counter$count = 94049;
	#10 counter$count = 94050;
	#10 counter$count = 94051;
	#10 counter$count = 94052;
	#10 counter$count = 94053;
	#10 counter$count = 94054;
	#10 counter$count = 94055;
	#10 counter$count = 94056;
	#10 counter$count = 94057;
	#10 counter$count = 94058;
	#10 counter$count = 94059;
	#10 counter$count = 94060;
	#10 counter$count = 94061;
	#10 counter$count = 94062;
	#10 counter$count = 94063;
	#10 counter$count = 94064;
	#10 counter$count = 94065;
	#10 counter$count = 94066;
	#10 counter$count = 94067;
	#10 counter$count = 94068;
	#10 counter$count = 94069;
	#10 counter$count = 94070;
	#10 counter$count = 94071;
	#10 counter$count = 94072;
	#10 counter$count = 94073;
	#10 counter$count = 94074;
	#10 counter$count = 94075;
	#10 counter$count = 94076;
	#10 counter$count = 94077;
	#10 counter$count = 94078;
	#10 counter$count = 94079;
	#10 counter$count = 94080;
	#10 counter$count = 94081;
	#10 counter$count = 94082;
	#10 counter$count = 94083;
	#10 counter$count = 94084;
	#10 counter$count = 94085;
	#10 counter$count = 94086;
	#10 counter$count = 94087;
	#10 counter$count = 94088;
	#10 counter$count = 94089;
	#10 counter$count = 94090;
	#10 counter$count = 94091;
	#10 counter$count = 94092;
	#10 counter$count = 94093;
	#10 counter$count = 94094;
	#10 counter$count = 94095;
	#10 counter$count = 94096;
	#10 counter$count = 94097;
	#10 counter$count = 94098;
	#10 counter$count = 94099;
	#10 counter$count = 94100;
	#10 counter$count = 94101;
	#10 counter$count = 94102;
	#10 counter$count = 94103;
	#10 counter$count = 94104;
	#10 counter$count = 94105;
	#10 counter$count = 94106;
	#10 counter$count = 94107;
	#10 counter$count = 94108;
	#10 counter$count = 94109;
	#10 counter$count = 94110;
	#10 counter$count = 94111;
	#10 counter$count = 94112;
	#10 counter$count = 94113;
	#10 counter$count = 94114;
	#10 counter$count = 94115;
	#10 counter$count = 94116;
	#10 counter$count = 94117;
	#10 counter$count = 94118;
	#10 counter$count = 94119;
	#10 counter$count = 94120;
	#10 counter$count = 94121;
	#10 counter$count = 94122;
	#10 counter$count = 94123;
	#10 counter$count = 94124;
	#10 counter$count = 94125;
	#10 counter$count = 94126;
	#10 counter$count = 94127;
	#10 counter$count = 94128;
	#10 counter$count = 94129;
	#10 counter$count = 94130;
	#10 counter$count = 94131;
	#10 counter$count = 94132;
	#10 counter$count = 94133;
	#10 counter$count = 94134;
	#10 counter$count = 94135;
	#10 counter$count = 94136;
	#10 counter$count = 94137;
	#10 counter$count = 94138;
	#10 counter$count = 94139;
	#10 counter$count = 94140;
	#10 counter$count = 94141;
	#10 counter$count = 94142;
	#10 counter$count = 94143;
	#10 counter$count = 94144;
	#10 counter$count = 94145;
	#10 counter$count = 94146;
	#10 counter$count = 94147;
	#10 counter$count = 94148;
	#10 counter$count = 94149;
	#10 counter$count = 94150;
	#10 counter$count = 94151;
	#10 counter$count = 94152;
	#10 counter$count = 94153;
	#10 counter$count = 94154;
	#10 counter$count = 94155;
	#10 counter$count = 94156;
	#10 counter$count = 94157;
	#10 counter$count = 94158;
	#10 counter$count = 94159;
	#10 counter$count = 94160;
	#10 counter$count = 94161;
	#10 counter$count = 94162;
	#10 counter$count = 94163;
	#10 counter$count = 94164;
	#10 counter$count = 94165;
	#10 counter$count = 94166;
	#10 counter$count = 94167;
	#10 counter$count = 94168;
	#10 counter$count = 94169;
	#10 counter$count = 94170;
	#10 counter$count = 94171;
	#10 counter$count = 94172;
	#10 counter$count = 94173;
	#10 counter$count = 94174;
	#10 counter$count = 94175;
	#10 counter$count = 94176;
	#10 counter$count = 94177;
	#10 counter$count = 94178;
	#10 counter$count = 94179;
	#10 counter$count = 94180;
	#10 counter$count = 94181;
	#10 counter$count = 94182;
	#10 counter$count = 94183;
	#10 counter$count = 94184;
	#10 counter$count = 94185;
	#10 counter$count = 94186;
	#10 counter$count = 94187;
	#10 counter$count = 94188;
	#10 counter$count = 94189;
	#10 counter$count = 94190;
	#10 counter$count = 94191;
	#10 counter$count = 94192;
	#10 counter$count = 94193;
	#10 counter$count = 94194;
	#10 counter$count = 94195;
	#10 counter$count = 94196;
	#10 counter$count = 94197;
	#10 counter$count = 94198;
	#10 counter$count = 94199;
	#10 counter$count = 94200;
	#10 counter$count = 94201;
	#10 counter$count = 94202;
	#10 counter$count = 94203;
	#10 counter$count = 94204;
	#10 counter$count = 94205;
	#10 counter$count = 94206;
	#10 counter$count = 94207;
	#10 counter$count = 94208;
	#10 counter$count = 94209;
	#10 counter$count = 94210;
	#10 counter$count = 94211;
	#10 counter$count = 94212;
	#10 counter$count = 94213;
	#10 counter$count = 94214;
	#10 counter$count = 94215;
	#10 counter$count = 94216;
	#10 counter$count = 94217;
	#10 counter$count = 94218;
	#10 counter$count = 94219;
	#10 counter$count = 94220;
	#10 counter$count = 94221;
	#10 counter$count = 94222;
	#10 counter$count = 94223;
	#10 counter$count = 94224;
	#10 counter$count = 94225;
	#10 counter$count = 94226;
	#10 counter$count = 94227;
	#10 counter$count = 94228;
	#10 counter$count = 94229;
	#10 counter$count = 94230;
	#10 counter$count = 94231;
	#10 counter$count = 94232;
	#10 counter$count = 94233;
	#10 counter$count = 94234;
	#10 counter$count = 94235;
	#10 counter$count = 94236;
	#10 counter$count = 94237;
	#10 counter$count = 94238;
	#10 counter$count = 94239;
	#10 counter$count = 94240;
	#10 counter$count = 94241;
	#10 counter$count = 94242;
	#10 counter$count = 94243;
	#10 counter$count = 94244;
	#10 counter$count = 94245;
	#10 counter$count = 94246;
	#10 counter$count = 94247;
	#10 counter$count = 94248;
	#10 counter$count = 94249;
	#10 counter$count = 94250;
	#10 counter$count = 94251;
	#10 counter$count = 94252;
	#10 counter$count = 94253;
	#10 counter$count = 94254;
	#10 counter$count = 94255;
	#10 counter$count = 94256;
	#10 counter$count = 94257;
	#10 counter$count = 94258;
	#10 counter$count = 94259;
	#10 counter$count = 94260;
	#10 counter$count = 94261;
	#10 counter$count = 94262;
	#10 counter$count = 94263;
	#10 counter$count = 94264;
	#10 counter$count = 94265;
	#10 counter$count = 94266;
	#10 counter$count = 94267;
	#10 counter$count = 94268;
	#10 counter$count = 94269;
	#10 counter$count = 94270;
	#10 counter$count = 94271;
	#10 counter$count = 94272;
	#10 counter$count = 94273;
	#10 counter$count = 94274;
	#10 counter$count = 94275;
	#10 counter$count = 94276;
	#10 counter$count = 94277;
	#10 counter$count = 94278;
	#10 counter$count = 94279;
	#10 counter$count = 94280;
	#10 counter$count = 94281;
	#10 counter$count = 94282;
	#10 counter$count = 94283;
	#10 counter$count = 94284;
	#10 counter$count = 94285;
	#10 counter$count = 94286;
	#10 counter$count = 94287;
	#10 counter$count = 94288;
	#10 counter$count = 94289;
	#10 counter$count = 94290;
	#10 counter$count = 94291;
	#10 counter$count = 94292;
	#10 counter$count = 94293;
	#10 counter$count = 94294;
	#10 counter$count = 94295;
	#10 counter$count = 94296;
	#10 counter$count = 94297;
	#10 counter$count = 94298;
	#10 counter$count = 94299;
	#10 counter$count = 94300;
	#10 counter$count = 94301;
	#10 counter$count = 94302;
	#10 counter$count = 94303;
	#10 counter$count = 94304;
	#10 counter$count = 94305;
	#10 counter$count = 94306;
	#10 counter$count = 94307;
	#10 counter$count = 94308;
	#10 counter$count = 94309;
	#10 counter$count = 94310;
	#10 counter$count = 94311;
	#10 counter$count = 94312;
	#10 counter$count = 94313;
	#10 counter$count = 94314;
	#10 counter$count = 94315;
	#10 counter$count = 94316;
	#10 counter$count = 94317;
	#10 counter$count = 94318;
	#10 counter$count = 94319;
	#10 counter$count = 94320;
	#10 counter$count = 94321;
	#10 counter$count = 94322;
	#10 counter$count = 94323;
	#10 counter$count = 94324;
	#10 counter$count = 94325;
	#10 counter$count = 94326;
	#10 counter$count = 94327;
	#10 counter$count = 94328;
	#10 counter$count = 94329;
	#10 counter$count = 94330;
	#10 counter$count = 94331;
	#10 counter$count = 94332;
	#10 counter$count = 94333;
	#10 counter$count = 94334;
	#10 counter$count = 94335;
	#10 counter$count = 94336;
	#10 counter$count = 94337;
	#10 counter$count = 94338;
	#10 counter$count = 94339;
	#10 counter$count = 94340;
	#10 counter$count = 94341;
	#10 counter$count = 94342;
	#10 counter$count = 94343;
	#10 counter$count = 94344;
	#10 counter$count = 94345;
	#10 counter$count = 94346;
	#10 counter$count = 94347;
	#10 counter$count = 94348;
	#10 counter$count = 94349;
	#10 counter$count = 94350;
	#10 counter$count = 94351;
	#10 counter$count = 94352;
	#10 counter$count = 94353;
	#10 counter$count = 94354;
	#10 counter$count = 94355;
	#10 counter$count = 94356;
	#10 counter$count = 94357;
	#10 counter$count = 94358;
	#10 counter$count = 94359;
	#10 counter$count = 94360;
	#10 counter$count = 94361;
	#10 counter$count = 94362;
	#10 counter$count = 94363;
	#10 counter$count = 94364;
	#10 counter$count = 94365;
	#10 counter$count = 94366;
	#10 counter$count = 94367;
	#10 counter$count = 94368;
	#10 counter$count = 94369;
	#10 counter$count = 94370;
	#10 counter$count = 94371;
	#10 counter$count = 94372;
	#10 counter$count = 94373;
	#10 counter$count = 94374;
	#10 counter$count = 94375;
	#10 counter$count = 94376;
	#10 counter$count = 94377;
	#10 counter$count = 94378;
	#10 counter$count = 94379;
	#10 counter$count = 94380;
	#10 counter$count = 94381;
	#10 counter$count = 94382;
	#10 counter$count = 94383;
	#10 counter$count = 94384;
	#10 counter$count = 94385;
	#10 counter$count = 94386;
	#10 counter$count = 94387;
	#10 counter$count = 94388;
	#10 counter$count = 94389;
	#10 counter$count = 94390;
	#10 counter$count = 94391;
	#10 counter$count = 94392;
	#10 counter$count = 94393;
	#10 counter$count = 94394;
	#10 counter$count = 94395;
	#10 counter$count = 94396;
	#10 counter$count = 94397;
	#10 counter$count = 94398;
	#10 counter$count = 94399;
	#10 counter$count = 94400;
	#10 counter$count = 94401;
	#10 counter$count = 94402;
	#10 counter$count = 94403;
	#10 counter$count = 94404;
	#10 counter$count = 94405;
	#10 counter$count = 94406;
	#10 counter$count = 94407;
	#10 counter$count = 94408;
	#10 counter$count = 94409;
	#10 counter$count = 94410;
	#10 counter$count = 94411;
	#10 counter$count = 94412;
	#10 counter$count = 94413;
	#10 counter$count = 94414;
	#10 counter$count = 94415;
	#10 counter$count = 94416;
	#10 counter$count = 94417;
	#10 counter$count = 94418;
	#10 counter$count = 94419;
	#10 counter$count = 94420;
	#10 counter$count = 94421;
	#10 counter$count = 94422;
	#10 counter$count = 94423;
	#10 counter$count = 94424;
	#10 counter$count = 94425;
	#10 counter$count = 94426;
	#10 counter$count = 94427;
	#10 counter$count = 94428;
	#10 counter$count = 94429;
	#10 counter$count = 94430;
	#10 counter$count = 94431;
	#10 counter$count = 94432;
	#10 counter$count = 94433;
	#10 counter$count = 94434;
	#10 counter$count = 94435;
	#10 counter$count = 94436;
	#10 counter$count = 94437;
	#10 counter$count = 94438;
	#10 counter$count = 94439;
	#10 counter$count = 94440;
	#10 counter$count = 94441;
	#10 counter$count = 94442;
	#10 counter$count = 94443;
	#10 counter$count = 94444;
	#10 counter$count = 94445;
	#10 counter$count = 94446;
	#10 counter$count = 94447;
	#10 counter$count = 94448;
	#10 counter$count = 94449;
	#10 counter$count = 94450;
	#10 counter$count = 94451;
	#10 counter$count = 94452;
	#10 counter$count = 94453;
	#10 counter$count = 94454;
	#10 counter$count = 94455;
	#10 counter$count = 94456;
	#10 counter$count = 94457;
	#10 counter$count = 94458;
	#10 counter$count = 94459;
	#10 counter$count = 94460;
	#10 counter$count = 94461;
	#10 counter$count = 94462;
	#10 counter$count = 94463;
	#10 counter$count = 94464;
	#10 counter$count = 94465;
	#10 counter$count = 94466;
	#10 counter$count = 94467;
	#10 counter$count = 94468;
	#10 counter$count = 94469;
	#10 counter$count = 94470;
	#10 counter$count = 94471;
	#10 counter$count = 94472;
	#10 counter$count = 94473;
	#10 counter$count = 94474;
	#10 counter$count = 94475;
	#10 counter$count = 94476;
	#10 counter$count = 94477;
	#10 counter$count = 94478;
	#10 counter$count = 94479;
	#10 counter$count = 94480;
	#10 counter$count = 94481;
	#10 counter$count = 94482;
	#10 counter$count = 94483;
	#10 counter$count = 94484;
	#10 counter$count = 94485;
	#10 counter$count = 94486;
	#10 counter$count = 94487;
	#10 counter$count = 94488;
	#10 counter$count = 94489;
	#10 counter$count = 94490;
	#10 counter$count = 94491;
	#10 counter$count = 94492;
	#10 counter$count = 94493;
	#10 counter$count = 94494;
	#10 counter$count = 94495;
	#10 counter$count = 94496;
	#10 counter$count = 94497;
	#10 counter$count = 94498;
	#10 counter$count = 94499;
	#10 counter$count = 94500;
	#10 counter$count = 94501;
	#10 counter$count = 94502;
	#10 counter$count = 94503;
	#10 counter$count = 94504;
	#10 counter$count = 94505;
	#10 counter$count = 94506;
	#10 counter$count = 94507;
	#10 counter$count = 94508;
	#10 counter$count = 94509;
	#10 counter$count = 94510;
	#10 counter$count = 94511;
	#10 counter$count = 94512;
	#10 counter$count = 94513;
	#10 counter$count = 94514;
	#10 counter$count = 94515;
	#10 counter$count = 94516;
	#10 counter$count = 94517;
	#10 counter$count = 94518;
	#10 counter$count = 94519;
	#10 counter$count = 94520;
	#10 counter$count = 94521;
	#10 counter$count = 94522;
	#10 counter$count = 94523;
	#10 counter$count = 94524;
	#10 counter$count = 94525;
	#10 counter$count = 94526;
	#10 counter$count = 94527;
	#10 counter$count = 94528;
	#10 counter$count = 94529;
	#10 counter$count = 94530;
	#10 counter$count = 94531;
	#10 counter$count = 94532;
	#10 counter$count = 94533;
	#10 counter$count = 94534;
	#10 counter$count = 94535;
	#10 counter$count = 94536;
	#10 counter$count = 94537;
	#10 counter$count = 94538;
	#10 counter$count = 94539;
	#10 counter$count = 94540;
	#10 counter$count = 94541;
	#10 counter$count = 94542;
	#10 counter$count = 94543;
	#10 counter$count = 94544;
	#10 counter$count = 94545;
	#10 counter$count = 94546;
	#10 counter$count = 94547;
	#10 counter$count = 94548;
	#10 counter$count = 94549;
	#10 counter$count = 94550;
	#10 counter$count = 94551;
	#10 counter$count = 94552;
	#10 counter$count = 94553;
	#10 counter$count = 94554;
	#10 counter$count = 94555;
	#10 counter$count = 94556;
	#10 counter$count = 94557;
	#10 counter$count = 94558;
	#10 counter$count = 94559;
	#10 counter$count = 94560;
	#10 counter$count = 94561;
	#10 counter$count = 94562;
	#10 counter$count = 94563;
	#10 counter$count = 94564;
	#10 counter$count = 94565;
	#10 counter$count = 94566;
	#10 counter$count = 94567;
	#10 counter$count = 94568;
	#10 counter$count = 94569;
	#10 counter$count = 94570;
	#10 counter$count = 94571;
	#10 counter$count = 94572;
	#10 counter$count = 94573;
	#10 counter$count = 94574;
	#10 counter$count = 94575;
	#10 counter$count = 94576;
	#10 counter$count = 94577;
	#10 counter$count = 94578;
	#10 counter$count = 94579;
	#10 counter$count = 94580;
	#10 counter$count = 94581;
	#10 counter$count = 94582;
	#10 counter$count = 94583;
	#10 counter$count = 94584;
	#10 counter$count = 94585;
	#10 counter$count = 94586;
	#10 counter$count = 94587;
	#10 counter$count = 94588;
	#10 counter$count = 94589;
	#10 counter$count = 94590;
	#10 counter$count = 94591;
	#10 counter$count = 94592;
	#10 counter$count = 94593;
	#10 counter$count = 94594;
	#10 counter$count = 94595;
	#10 counter$count = 94596;
	#10 counter$count = 94597;
	#10 counter$count = 94598;
	#10 counter$count = 94599;
	#10 counter$count = 94600;
	#10 counter$count = 94601;
	#10 counter$count = 94602;
	#10 counter$count = 94603;
	#10 counter$count = 94604;
	#10 counter$count = 94605;
	#10 counter$count = 94606;
	#10 counter$count = 94607;
	#10 counter$count = 94608;
	#10 counter$count = 94609;
	#10 counter$count = 94610;
	#10 counter$count = 94611;
	#10 counter$count = 94612;
	#10 counter$count = 94613;
	#10 counter$count = 94614;
	#10 counter$count = 94615;
	#10 counter$count = 94616;
	#10 counter$count = 94617;
	#10 counter$count = 94618;
	#10 counter$count = 94619;
	#10 counter$count = 94620;
	#10 counter$count = 94621;
	#10 counter$count = 94622;
	#10 counter$count = 94623;
	#10 counter$count = 94624;
	#10 counter$count = 94625;
	#10 counter$count = 94626;
	#10 counter$count = 94627;
	#10 counter$count = 94628;
	#10 counter$count = 94629;
	#10 counter$count = 94630;
	#10 counter$count = 94631;
	#10 counter$count = 94632;
	#10 counter$count = 94633;
	#10 counter$count = 94634;
	#10 counter$count = 94635;
	#10 counter$count = 94636;
	#10 counter$count = 94637;
	#10 counter$count = 94638;
	#10 counter$count = 94639;
	#10 counter$count = 94640;
	#10 counter$count = 94641;
	#10 counter$count = 94642;
	#10 counter$count = 94643;
	#10 counter$count = 94644;
	#10 counter$count = 94645;
	#10 counter$count = 94646;
	#10 counter$count = 94647;
	#10 counter$count = 94648;
	#10 counter$count = 94649;
	#10 counter$count = 94650;
	#10 counter$count = 94651;
	#10 counter$count = 94652;
	#10 counter$count = 94653;
	#10 counter$count = 94654;
	#10 counter$count = 94655;
	#10 counter$count = 94656;
	#10 counter$count = 94657;
	#10 counter$count = 94658;
	#10 counter$count = 94659;
	#10 counter$count = 94660;
	#10 counter$count = 94661;
	#10 counter$count = 94662;
	#10 counter$count = 94663;
	#10 counter$count = 94664;
	#10 counter$count = 94665;
	#10 counter$count = 94666;
	#10 counter$count = 94667;
	#10 counter$count = 94668;
	#10 counter$count = 94669;
	#10 counter$count = 94670;
	#10 counter$count = 94671;
	#10 counter$count = 94672;
	#10 counter$count = 94673;
	#10 counter$count = 94674;
	#10 counter$count = 94675;
	#10 counter$count = 94676;
	#10 counter$count = 94677;
	#10 counter$count = 94678;
	#10 counter$count = 94679;
	#10 counter$count = 94680;
	#10 counter$count = 94681;
	#10 counter$count = 94682;
	#10 counter$count = 94683;
	#10 counter$count = 94684;
	#10 counter$count = 94685;
	#10 counter$count = 94686;
	#10 counter$count = 94687;
	#10 counter$count = 94688;
	#10 counter$count = 94689;
	#10 counter$count = 94690;
	#10 counter$count = 94691;
	#10 counter$count = 94692;
	#10 counter$count = 94693;
	#10 counter$count = 94694;
	#10 counter$count = 94695;
	#10 counter$count = 94696;
	#10 counter$count = 94697;
	#10 counter$count = 94698;
	#10 counter$count = 94699;
	#10 counter$count = 94700;
	#10 counter$count = 94701;
	#10 counter$count = 94702;
	#10 counter$count = 94703;
	#10 counter$count = 94704;
	#10 counter$count = 94705;
	#10 counter$count = 94706;
	#10 counter$count = 94707;
	#10 counter$count = 94708;
	#10 counter$count = 94709;
	#10 counter$count = 94710;
	#10 counter$count = 94711;
	#10 counter$count = 94712;
	#10 counter$count = 94713;
	#10 counter$count = 94714;
	#10 counter$count = 94715;
	#10 counter$count = 94716;
	#10 counter$count = 94717;
	#10 counter$count = 94718;
	#10 counter$count = 94719;
	#10 counter$count = 94720;
	#10 counter$count = 94721;
	#10 counter$count = 94722;
	#10 counter$count = 94723;
	#10 counter$count = 94724;
	#10 counter$count = 94725;
	#10 counter$count = 94726;
	#10 counter$count = 94727;
	#10 counter$count = 94728;
	#10 counter$count = 94729;
	#10 counter$count = 94730;
	#10 counter$count = 94731;
	#10 counter$count = 94732;
	#10 counter$count = 94733;
	#10 counter$count = 94734;
	#10 counter$count = 94735;
	#10 counter$count = 94736;
	#10 counter$count = 94737;
	#10 counter$count = 94738;
	#10 counter$count = 94739;
	#10 counter$count = 94740;
	#10 counter$count = 94741;
	#10 counter$count = 94742;
	#10 counter$count = 94743;
	#10 counter$count = 94744;
	#10 counter$count = 94745;
	#10 counter$count = 94746;
	#10 counter$count = 94747;
	#10 counter$count = 94748;
	#10 counter$count = 94749;
	#10 counter$count = 94750;
	#10 counter$count = 94751;
	#10 counter$count = 94752;
	#10 counter$count = 94753;
	#10 counter$count = 94754;
	#10 counter$count = 94755;
	#10 counter$count = 94756;
	#10 counter$count = 94757;
	#10 counter$count = 94758;
	#10 counter$count = 94759;
	#10 counter$count = 94760;
	#10 counter$count = 94761;
	#10 counter$count = 94762;
	#10 counter$count = 94763;
	#10 counter$count = 94764;
	#10 counter$count = 94765;
	#10 counter$count = 94766;
	#10 counter$count = 94767;
	#10 counter$count = 94768;
	#10 counter$count = 94769;
	#10 counter$count = 94770;
	#10 counter$count = 94771;
	#10 counter$count = 94772;
	#10 counter$count = 94773;
	#10 counter$count = 94774;
	#10 counter$count = 94775;
	#10 counter$count = 94776;
	#10 counter$count = 94777;
	#10 counter$count = 94778;
	#10 counter$count = 94779;
	#10 counter$count = 94780;
	#10 counter$count = 94781;
	#10 counter$count = 94782;
	#10 counter$count = 94783;
	#10 counter$count = 94784;
	#10 counter$count = 94785;
	#10 counter$count = 94786;
	#10 counter$count = 94787;
	#10 counter$count = 94788;
	#10 counter$count = 94789;
	#10 counter$count = 94790;
	#10 counter$count = 94791;
	#10 counter$count = 94792;
	#10 counter$count = 94793;
	#10 counter$count = 94794;
	#10 counter$count = 94795;
	#10 counter$count = 94796;
	#10 counter$count = 94797;
	#10 counter$count = 94798;
	#10 counter$count = 94799;
	#10 counter$count = 94800;
	#10 counter$count = 94801;
	#10 counter$count = 94802;
	#10 counter$count = 94803;
	#10 counter$count = 94804;
	#10 counter$count = 94805;
	#10 counter$count = 94806;
	#10 counter$count = 94807;
	#10 counter$count = 94808;
	#10 counter$count = 94809;
	#10 counter$count = 94810;
	#10 counter$count = 94811;
	#10 counter$count = 94812;
	#10 counter$count = 94813;
	#10 counter$count = 94814;
	#10 counter$count = 94815;
	#10 counter$count = 94816;
	#10 counter$count = 94817;
	#10 counter$count = 94818;
	#10 counter$count = 94819;
	#10 counter$count = 94820;
	#10 counter$count = 94821;
	#10 counter$count = 94822;
	#10 counter$count = 94823;
	#10 counter$count = 94824;
	#10 counter$count = 94825;
	#10 counter$count = 94826;
	#10 counter$count = 94827;
	#10 counter$count = 94828;
	#10 counter$count = 94829;
	#10 counter$count = 94830;
	#10 counter$count = 94831;
	#10 counter$count = 94832;
	#10 counter$count = 94833;
	#10 counter$count = 94834;
	#10 counter$count = 94835;
	#10 counter$count = 94836;
	#10 counter$count = 94837;
	#10 counter$count = 94838;
	#10 counter$count = 94839;
	#10 counter$count = 94840;
	#10 counter$count = 94841;
	#10 counter$count = 94842;
	#10 counter$count = 94843;
	#10 counter$count = 94844;
	#10 counter$count = 94845;
	#10 counter$count = 94846;
	#10 counter$count = 94847;
	#10 counter$count = 94848;
	#10 counter$count = 94849;
	#10 counter$count = 94850;
	#10 counter$count = 94851;
	#10 counter$count = 94852;
	#10 counter$count = 94853;
	#10 counter$count = 94854;
	#10 counter$count = 94855;
	#10 counter$count = 94856;
	#10 counter$count = 94857;
	#10 counter$count = 94858;
	#10 counter$count = 94859;
	#10 counter$count = 94860;
	#10 counter$count = 94861;
	#10 counter$count = 94862;
	#10 counter$count = 94863;
	#10 counter$count = 94864;
	#10 counter$count = 94865;
	#10 counter$count = 94866;
	#10 counter$count = 94867;
	#10 counter$count = 94868;
	#10 counter$count = 94869;
	#10 counter$count = 94870;
	#10 counter$count = 94871;
	#10 counter$count = 94872;
	#10 counter$count = 94873;
	#10 counter$count = 94874;
	#10 counter$count = 94875;
	#10 counter$count = 94876;
	#10 counter$count = 94877;
	#10 counter$count = 94878;
	#10 counter$count = 94879;
	#10 counter$count = 94880;
	#10 counter$count = 94881;
	#10 counter$count = 94882;
	#10 counter$count = 94883;
	#10 counter$count = 94884;
	#10 counter$count = 94885;
	#10 counter$count = 94886;
	#10 counter$count = 94887;
	#10 counter$count = 94888;
	#10 counter$count = 94889;
	#10 counter$count = 94890;
	#10 counter$count = 94891;
	#10 counter$count = 94892;
	#10 counter$count = 94893;
	#10 counter$count = 94894;
	#10 counter$count = 94895;
	#10 counter$count = 94896;
	#10 counter$count = 94897;
	#10 counter$count = 94898;
	#10 counter$count = 94899;
	#10 counter$count = 94900;
	#10 counter$count = 94901;
	#10 counter$count = 94902;
	#10 counter$count = 94903;
	#10 counter$count = 94904;
	#10 counter$count = 94905;
	#10 counter$count = 94906;
	#10 counter$count = 94907;
	#10 counter$count = 94908;
	#10 counter$count = 94909;
	#10 counter$count = 94910;
	#10 counter$count = 94911;
	#10 counter$count = 94912;
	#10 counter$count = 94913;
	#10 counter$count = 94914;
	#10 counter$count = 94915;
	#10 counter$count = 94916;
	#10 counter$count = 94917;
	#10 counter$count = 94918;
	#10 counter$count = 94919;
	#10 counter$count = 94920;
	#10 counter$count = 94921;
	#10 counter$count = 94922;
	#10 counter$count = 94923;
	#10 counter$count = 94924;
	#10 counter$count = 94925;
	#10 counter$count = 94926;
	#10 counter$count = 94927;
	#10 counter$count = 94928;
	#10 counter$count = 94929;
	#10 counter$count = 94930;
	#10 counter$count = 94931;
	#10 counter$count = 94932;
	#10 counter$count = 94933;
	#10 counter$count = 94934;
	#10 counter$count = 94935;
	#10 counter$count = 94936;
	#10 counter$count = 94937;
	#10 counter$count = 94938;
	#10 counter$count = 94939;
	#10 counter$count = 94940;
	#10 counter$count = 94941;
	#10 counter$count = 94942;
	#10 counter$count = 94943;
	#10 counter$count = 94944;
	#10 counter$count = 94945;
	#10 counter$count = 94946;
	#10 counter$count = 94947;
	#10 counter$count = 94948;
	#10 counter$count = 94949;
	#10 counter$count = 94950;
	#10 counter$count = 94951;
	#10 counter$count = 94952;
	#10 counter$count = 94953;
	#10 counter$count = 94954;
	#10 counter$count = 94955;
	#10 counter$count = 94956;
	#10 counter$count = 94957;
	#10 counter$count = 94958;
	#10 counter$count = 94959;
	#10 counter$count = 94960;
	#10 counter$count = 94961;
	#10 counter$count = 94962;
	#10 counter$count = 94963;
	#10 counter$count = 94964;
	#10 counter$count = 94965;
	#10 counter$count = 94966;
	#10 counter$count = 94967;
	#10 counter$count = 94968;
	#10 counter$count = 94969;
	#10 counter$count = 94970;
	#10 counter$count = 94971;
	#10 counter$count = 94972;
	#10 counter$count = 94973;
	#10 counter$count = 94974;
	#10 counter$count = 94975;
	#10 counter$count = 94976;
	#10 counter$count = 94977;
	#10 counter$count = 94978;
	#10 counter$count = 94979;
	#10 counter$count = 94980;
	#10 counter$count = 94981;
	#10 counter$count = 94982;
	#10 counter$count = 94983;
	#10 counter$count = 94984;
	#10 counter$count = 94985;
	#10 counter$count = 94986;
	#10 counter$count = 94987;
	#10 counter$count = 94988;
	#10 counter$count = 94989;
	#10 counter$count = 94990;
	#10 counter$count = 94991;
	#10 counter$count = 94992;
	#10 counter$count = 94993;
	#10 counter$count = 94994;
	#10 counter$count = 94995;
	#10 counter$count = 94996;
	#10 counter$count = 94997;
	#10 counter$count = 94998;
	#10 counter$count = 94999;
	#10 counter$count = 95000;
	#10 counter$count = 95001;
	#10 counter$count = 95002;
	#10 counter$count = 95003;
	#10 counter$count = 95004;
	#10 counter$count = 95005;
	#10 counter$count = 95006;
	#10 counter$count = 95007;
	#10 counter$count = 95008;
	#10 counter$count = 95009;
	#10 counter$count = 95010;
	#10 counter$count = 95011;
	#10 counter$count = 95012;
	#10 counter$count = 95013;
	#10 counter$count = 95014;
	#10 counter$count = 95015;
	#10 counter$count = 95016;
	#10 counter$count = 95017;
	#10 counter$count = 95018;
	#10 counter$count = 95019;
	#10 counter$count = 95020;
	#10 counter$count = 95021;
	#10 counter$count = 95022;
	#10 counter$count = 95023;
	#10 counter$count = 95024;
	#10 counter$count = 95025;
	#10 counter$count = 95026;
	#10 counter$count = 95027;
	#10 counter$count = 95028;
	#10 counter$count = 95029;
	#10 counter$count = 95030;
	#10 counter$count = 95031;
	#10 counter$count = 95032;
	#10 counter$count = 95033;
	#10 counter$count = 95034;
	#10 counter$count = 95035;
	#10 counter$count = 95036;
	#10 counter$count = 95037;
	#10 counter$count = 95038;
	#10 counter$count = 95039;
	#10 counter$count = 95040;
	#10 counter$count = 95041;
	#10 counter$count = 95042;
	#10 counter$count = 95043;
	#10 counter$count = 95044;
	#10 counter$count = 95045;
	#10 counter$count = 95046;
	#10 counter$count = 95047;
	#10 counter$count = 95048;
	#10 counter$count = 95049;
	#10 counter$count = 95050;
	#10 counter$count = 95051;
	#10 counter$count = 95052;
	#10 counter$count = 95053;
	#10 counter$count = 95054;
	#10 counter$count = 95055;
	#10 counter$count = 95056;
	#10 counter$count = 95057;
	#10 counter$count = 95058;
	#10 counter$count = 95059;
	#10 counter$count = 95060;
	#10 counter$count = 95061;
	#10 counter$count = 95062;
	#10 counter$count = 95063;
	#10 counter$count = 95064;
	#10 counter$count = 95065;
	#10 counter$count = 95066;
	#10 counter$count = 95067;
	#10 counter$count = 95068;
	#10 counter$count = 95069;
	#10 counter$count = 95070;
	#10 counter$count = 95071;
	#10 counter$count = 95072;
	#10 counter$count = 95073;
	#10 counter$count = 95074;
	#10 counter$count = 95075;
	#10 counter$count = 95076;
	#10 counter$count = 95077;
	#10 counter$count = 95078;
	#10 counter$count = 95079;
	#10 counter$count = 95080;
	#10 counter$count = 95081;
	#10 counter$count = 95082;
	#10 counter$count = 95083;
	#10 counter$count = 95084;
	#10 counter$count = 95085;
	#10 counter$count = 95086;
	#10 counter$count = 95087;
	#10 counter$count = 95088;
	#10 counter$count = 95089;
	#10 counter$count = 95090;
	#10 counter$count = 95091;
	#10 counter$count = 95092;
	#10 counter$count = 95093;
	#10 counter$count = 95094;
	#10 counter$count = 95095;
	#10 counter$count = 95096;
	#10 counter$count = 95097;
	#10 counter$count = 95098;
	#10 counter$count = 95099;
	#10 counter$count = 95100;
	#10 counter$count = 95101;
	#10 counter$count = 95102;
	#10 counter$count = 95103;
	#10 counter$count = 95104;
	#10 counter$count = 95105;
	#10 counter$count = 95106;
	#10 counter$count = 95107;
	#10 counter$count = 95108;
	#10 counter$count = 95109;
	#10 counter$count = 95110;
	#10 counter$count = 95111;
	#10 counter$count = 95112;
	#10 counter$count = 95113;
	#10 counter$count = 95114;
	#10 counter$count = 95115;
	#10 counter$count = 95116;
	#10 counter$count = 95117;
	#10 counter$count = 95118;
	#10 counter$count = 95119;
	#10 counter$count = 95120;
	#10 counter$count = 95121;
	#10 counter$count = 95122;
	#10 counter$count = 95123;
	#10 counter$count = 95124;
	#10 counter$count = 95125;
	#10 counter$count = 95126;
	#10 counter$count = 95127;
	#10 counter$count = 95128;
	#10 counter$count = 95129;
	#10 counter$count = 95130;
	#10 counter$count = 95131;
	#10 counter$count = 95132;
	#10 counter$count = 95133;
	#10 counter$count = 95134;
	#10 counter$count = 95135;
	#10 counter$count = 95136;
	#10 counter$count = 95137;
	#10 counter$count = 95138;
	#10 counter$count = 95139;
	#10 counter$count = 95140;
	#10 counter$count = 95141;
	#10 counter$count = 95142;
	#10 counter$count = 95143;
	#10 counter$count = 95144;
	#10 counter$count = 95145;
	#10 counter$count = 95146;
	#10 counter$count = 95147;
	#10 counter$count = 95148;
	#10 counter$count = 95149;
	#10 counter$count = 95150;
	#10 counter$count = 95151;
	#10 counter$count = 95152;
	#10 counter$count = 95153;
	#10 counter$count = 95154;
	#10 counter$count = 95155;
	#10 counter$count = 95156;
	#10 counter$count = 95157;
	#10 counter$count = 95158;
	#10 counter$count = 95159;
	#10 counter$count = 95160;
	#10 counter$count = 95161;
	#10 counter$count = 95162;
	#10 counter$count = 95163;
	#10 counter$count = 95164;
	#10 counter$count = 95165;
	#10 counter$count = 95166;
	#10 counter$count = 95167;
	#10 counter$count = 95168;
	#10 counter$count = 95169;
	#10 counter$count = 95170;
	#10 counter$count = 95171;
	#10 counter$count = 95172;
	#10 counter$count = 95173;
	#10 counter$count = 95174;
	#10 counter$count = 95175;
	#10 counter$count = 95176;
	#10 counter$count = 95177;
	#10 counter$count = 95178;
	#10 counter$count = 95179;
	#10 counter$count = 95180;
	#10 counter$count = 95181;
	#10 counter$count = 95182;
	#10 counter$count = 95183;
	#10 counter$count = 95184;
	#10 counter$count = 95185;
	#10 counter$count = 95186;
	#10 counter$count = 95187;
	#10 counter$count = 95188;
	#10 counter$count = 95189;
	#10 counter$count = 95190;
	#10 counter$count = 95191;
	#10 counter$count = 95192;
	#10 counter$count = 95193;
	#10 counter$count = 95194;
	#10 counter$count = 95195;
	#10 counter$count = 95196;
	#10 counter$count = 95197;
	#10 counter$count = 95198;
	#10 counter$count = 95199;
	#10 counter$count = 95200;
	#10 counter$count = 95201;
	#10 counter$count = 95202;
	#10 counter$count = 95203;
	#10 counter$count = 95204;
	#10 counter$count = 95205;
	#10 counter$count = 95206;
	#10 counter$count = 95207;
	#10 counter$count = 95208;
	#10 counter$count = 95209;
	#10 counter$count = 95210;
	#10 counter$count = 95211;
	#10 counter$count = 95212;
	#10 counter$count = 95213;
	#10 counter$count = 95214;
	#10 counter$count = 95215;
	#10 counter$count = 95216;
	#10 counter$count = 95217;
	#10 counter$count = 95218;
	#10 counter$count = 95219;
	#10 counter$count = 95220;
	#10 counter$count = 95221;
	#10 counter$count = 95222;
	#10 counter$count = 95223;
	#10 counter$count = 95224;
	#10 counter$count = 95225;
	#10 counter$count = 95226;
	#10 counter$count = 95227;
	#10 counter$count = 95228;
	#10 counter$count = 95229;
	#10 counter$count = 95230;
	#10 counter$count = 95231;
	#10 counter$count = 95232;
	#10 counter$count = 95233;
	#10 counter$count = 95234;
	#10 counter$count = 95235;
	#10 counter$count = 95236;
	#10 counter$count = 95237;
	#10 counter$count = 95238;
	#10 counter$count = 95239;
	#10 counter$count = 95240;
	#10 counter$count = 95241;
	#10 counter$count = 95242;
	#10 counter$count = 95243;
	#10 counter$count = 95244;
	#10 counter$count = 95245;
	#10 counter$count = 95246;
	#10 counter$count = 95247;
	#10 counter$count = 95248;
	#10 counter$count = 95249;
	#10 counter$count = 95250;
	#10 counter$count = 95251;
	#10 counter$count = 95252;
	#10 counter$count = 95253;
	#10 counter$count = 95254;
	#10 counter$count = 95255;
	#10 counter$count = 95256;
	#10 counter$count = 95257;
	#10 counter$count = 95258;
	#10 counter$count = 95259;
	#10 counter$count = 95260;
	#10 counter$count = 95261;
	#10 counter$count = 95262;
	#10 counter$count = 95263;
	#10 counter$count = 95264;
	#10 counter$count = 95265;
	#10 counter$count = 95266;
	#10 counter$count = 95267;
	#10 counter$count = 95268;
	#10 counter$count = 95269;
	#10 counter$count = 95270;
	#10 counter$count = 95271;
	#10 counter$count = 95272;
	#10 counter$count = 95273;
	#10 counter$count = 95274;
	#10 counter$count = 95275;
	#10 counter$count = 95276;
	#10 counter$count = 95277;
	#10 counter$count = 95278;
	#10 counter$count = 95279;
	#10 counter$count = 95280;
	#10 counter$count = 95281;
	#10 counter$count = 95282;
	#10 counter$count = 95283;
	#10 counter$count = 95284;
	#10 counter$count = 95285;
	#10 counter$count = 95286;
	#10 counter$count = 95287;
	#10 counter$count = 95288;
	#10 counter$count = 95289;
	#10 counter$count = 95290;
	#10 counter$count = 95291;
	#10 counter$count = 95292;
	#10 counter$count = 95293;
	#10 counter$count = 95294;
	#10 counter$count = 95295;
	#10 counter$count = 95296;
	#10 counter$count = 95297;
	#10 counter$count = 95298;
	#10 counter$count = 95299;
	#10 counter$count = 95300;
	#10 counter$count = 95301;
	#10 counter$count = 95302;
	#10 counter$count = 95303;
	#10 counter$count = 95304;
	#10 counter$count = 95305;
	#10 counter$count = 95306;
	#10 counter$count = 95307;
	#10 counter$count = 95308;
	#10 counter$count = 95309;
	#10 counter$count = 95310;
	#10 counter$count = 95311;
	#10 counter$count = 95312;
	#10 counter$count = 95313;
	#10 counter$count = 95314;
	#10 counter$count = 95315;
	#10 counter$count = 95316;
	#10 counter$count = 95317;
	#10 counter$count = 95318;
	#10 counter$count = 95319;
	#10 counter$count = 95320;
	#10 counter$count = 95321;
	#10 counter$count = 95322;
	#10 counter$count = 95323;
	#10 counter$count = 95324;
	#10 counter$count = 95325;
	#10 counter$count = 95326;
	#10 counter$count = 95327;
	#10 counter$count = 95328;
	#10 counter$count = 95329;
	#10 counter$count = 95330;
	#10 counter$count = 95331;
	#10 counter$count = 95332;
	#10 counter$count = 95333;
	#10 counter$count = 95334;
	#10 counter$count = 95335;
	#10 counter$count = 95336;
	#10 counter$count = 95337;
	#10 counter$count = 95338;
	#10 counter$count = 95339;
	#10 counter$count = 95340;
	#10 counter$count = 95341;
	#10 counter$count = 95342;
	#10 counter$count = 95343;
	#10 counter$count = 95344;
	#10 counter$count = 95345;
	#10 counter$count = 95346;
	#10 counter$count = 95347;
	#10 counter$count = 95348;
	#10 counter$count = 95349;
	#10 counter$count = 95350;
	#10 counter$count = 95351;
	#10 counter$count = 95352;
	#10 counter$count = 95353;
	#10 counter$count = 95354;
	#10 counter$count = 95355;
	#10 counter$count = 95356;
	#10 counter$count = 95357;
	#10 counter$count = 95358;
	#10 counter$count = 95359;
	#10 counter$count = 95360;
	#10 counter$count = 95361;
	#10 counter$count = 95362;
	#10 counter$count = 95363;
	#10 counter$count = 95364;
	#10 counter$count = 95365;
	#10 counter$count = 95366;
	#10 counter$count = 95367;
	#10 counter$count = 95368;
	#10 counter$count = 95369;
	#10 counter$count = 95370;
	#10 counter$count = 95371;
	#10 counter$count = 95372;
	#10 counter$count = 95373;
	#10 counter$count = 95374;
	#10 counter$count = 95375;
	#10 counter$count = 95376;
	#10 counter$count = 95377;
	#10 counter$count = 95378;
	#10 counter$count = 95379;
	#10 counter$count = 95380;
	#10 counter$count = 95381;
	#10 counter$count = 95382;
	#10 counter$count = 95383;
	#10 counter$count = 95384;
	#10 counter$count = 95385;
	#10 counter$count = 95386;
	#10 counter$count = 95387;
	#10 counter$count = 95388;
	#10 counter$count = 95389;
	#10 counter$count = 95390;
	#10 counter$count = 95391;
	#10 counter$count = 95392;
	#10 counter$count = 95393;
	#10 counter$count = 95394;
	#10 counter$count = 95395;
	#10 counter$count = 95396;
	#10 counter$count = 95397;
	#10 counter$count = 95398;
	#10 counter$count = 95399;
	#10 counter$count = 95400;
	#10 counter$count = 95401;
	#10 counter$count = 95402;
	#10 counter$count = 95403;
	#10 counter$count = 95404;
	#10 counter$count = 95405;
	#10 counter$count = 95406;
	#10 counter$count = 95407;
	#10 counter$count = 95408;
	#10 counter$count = 95409;
	#10 counter$count = 95410;
	#10 counter$count = 95411;
	#10 counter$count = 95412;
	#10 counter$count = 95413;
	#10 counter$count = 95414;
	#10 counter$count = 95415;
	#10 counter$count = 95416;
	#10 counter$count = 95417;
	#10 counter$count = 95418;
	#10 counter$count = 95419;
	#10 counter$count = 95420;
	#10 counter$count = 95421;
	#10 counter$count = 95422;
	#10 counter$count = 95423;
	#10 counter$count = 95424;
	#10 counter$count = 95425;
	#10 counter$count = 95426;
	#10 counter$count = 95427;
	#10 counter$count = 95428;
	#10 counter$count = 95429;
	#10 counter$count = 95430;
	#10 counter$count = 95431;
	#10 counter$count = 95432;
	#10 counter$count = 95433;
	#10 counter$count = 95434;
	#10 counter$count = 95435;
	#10 counter$count = 95436;
	#10 counter$count = 95437;
	#10 counter$count = 95438;
	#10 counter$count = 95439;
	#10 counter$count = 95440;
	#10 counter$count = 95441;
	#10 counter$count = 95442;
	#10 counter$count = 95443;
	#10 counter$count = 95444;
	#10 counter$count = 95445;
	#10 counter$count = 95446;
	#10 counter$count = 95447;
	#10 counter$count = 95448;
	#10 counter$count = 95449;
	#10 counter$count = 95450;
	#10 counter$count = 95451;
	#10 counter$count = 95452;
	#10 counter$count = 95453;
	#10 counter$count = 95454;
	#10 counter$count = 95455;
	#10 counter$count = 95456;
	#10 counter$count = 95457;
	#10 counter$count = 95458;
	#10 counter$count = 95459;
	#10 counter$count = 95460;
	#10 counter$count = 95461;
	#10 counter$count = 95462;
	#10 counter$count = 95463;
	#10 counter$count = 95464;
	#10 counter$count = 95465;
	#10 counter$count = 95466;
	#10 counter$count = 95467;
	#10 counter$count = 95468;
	#10 counter$count = 95469;
	#10 counter$count = 95470;
	#10 counter$count = 95471;
	#10 counter$count = 95472;
	#10 counter$count = 95473;
	#10 counter$count = 95474;
	#10 counter$count = 95475;
	#10 counter$count = 95476;
	#10 counter$count = 95477;
	#10 counter$count = 95478;
	#10 counter$count = 95479;
	#10 counter$count = 95480;
	#10 counter$count = 95481;
	#10 counter$count = 95482;
	#10 counter$count = 95483;
	#10 counter$count = 95484;
	#10 counter$count = 95485;
	#10 counter$count = 95486;
	#10 counter$count = 95487;
	#10 counter$count = 95488;
	#10 counter$count = 95489;
	#10 counter$count = 95490;
	#10 counter$count = 95491;
	#10 counter$count = 95492;
	#10 counter$count = 95493;
	#10 counter$count = 95494;
	#10 counter$count = 95495;
	#10 counter$count = 95496;
	#10 counter$count = 95497;
	#10 counter$count = 95498;
	#10 counter$count = 95499;
	#10 counter$count = 95500;
	#10 counter$count = 95501;
	#10 counter$count = 95502;
	#10 counter$count = 95503;
	#10 counter$count = 95504;
	#10 counter$count = 95505;
	#10 counter$count = 95506;
	#10 counter$count = 95507;
	#10 counter$count = 95508;
	#10 counter$count = 95509;
	#10 counter$count = 95510;
	#10 counter$count = 95511;
	#10 counter$count = 95512;
	#10 counter$count = 95513;
	#10 counter$count = 95514;
	#10 counter$count = 95515;
	#10 counter$count = 95516;
	#10 counter$count = 95517;
	#10 counter$count = 95518;
	#10 counter$count = 95519;
	#10 counter$count = 95520;
	#10 counter$count = 95521;
	#10 counter$count = 95522;
	#10 counter$count = 95523;
	#10 counter$count = 95524;
	#10 counter$count = 95525;
	#10 counter$count = 95526;
	#10 counter$count = 95527;
	#10 counter$count = 95528;
	#10 counter$count = 95529;
	#10 counter$count = 95530;
	#10 counter$count = 95531;
	#10 counter$count = 95532;
	#10 counter$count = 95533;
	#10 counter$count = 95534;
	#10 counter$count = 95535;
	#10 counter$count = 95536;
	#10 counter$count = 95537;
	#10 counter$count = 95538;
	#10 counter$count = 95539;
	#10 counter$count = 95540;
	#10 counter$count = 95541;
	#10 counter$count = 95542;
	#10 counter$count = 95543;
	#10 counter$count = 95544;
	#10 counter$count = 95545;
	#10 counter$count = 95546;
	#10 counter$count = 95547;
	#10 counter$count = 95548;
	#10 counter$count = 95549;
	#10 counter$count = 95550;
	#10 counter$count = 95551;
	#10 counter$count = 95552;
	#10 counter$count = 95553;
	#10 counter$count = 95554;
	#10 counter$count = 95555;
	#10 counter$count = 95556;
	#10 counter$count = 95557;
	#10 counter$count = 95558;
	#10 counter$count = 95559;
	#10 counter$count = 95560;
	#10 counter$count = 95561;
	#10 counter$count = 95562;
	#10 counter$count = 95563;
	#10 counter$count = 95564;
	#10 counter$count = 95565;
	#10 counter$count = 95566;
	#10 counter$count = 95567;
	#10 counter$count = 95568;
	#10 counter$count = 95569;
	#10 counter$count = 95570;
	#10 counter$count = 95571;
	#10 counter$count = 95572;
	#10 counter$count = 95573;
	#10 counter$count = 95574;
	#10 counter$count = 95575;
	#10 counter$count = 95576;
	#10 counter$count = 95577;
	#10 counter$count = 95578;
	#10 counter$count = 95579;
	#10 counter$count = 95580;
	#10 counter$count = 95581;
	#10 counter$count = 95582;
	#10 counter$count = 95583;
	#10 counter$count = 95584;
	#10 counter$count = 95585;
	#10 counter$count = 95586;
	#10 counter$count = 95587;
	#10 counter$count = 95588;
	#10 counter$count = 95589;
	#10 counter$count = 95590;
	#10 counter$count = 95591;
	#10 counter$count = 95592;
	#10 counter$count = 95593;
	#10 counter$count = 95594;
	#10 counter$count = 95595;
	#10 counter$count = 95596;
	#10 counter$count = 95597;
	#10 counter$count = 95598;
	#10 counter$count = 95599;
	#10 counter$count = 95600;
	#10 counter$count = 95601;
	#10 counter$count = 95602;
	#10 counter$count = 95603;
	#10 counter$count = 95604;
	#10 counter$count = 95605;
	#10 counter$count = 95606;
	#10 counter$count = 95607;
	#10 counter$count = 95608;
	#10 counter$count = 95609;
	#10 counter$count = 95610;
	#10 counter$count = 95611;
	#10 counter$count = 95612;
	#10 counter$count = 95613;
	#10 counter$count = 95614;
	#10 counter$count = 95615;
	#10 counter$count = 95616;
	#10 counter$count = 95617;
	#10 counter$count = 95618;
	#10 counter$count = 95619;
	#10 counter$count = 95620;
	#10 counter$count = 95621;
	#10 counter$count = 95622;
	#10 counter$count = 95623;
	#10 counter$count = 95624;
	#10 counter$count = 95625;
	#10 counter$count = 95626;
	#10 counter$count = 95627;
	#10 counter$count = 95628;
	#10 counter$count = 95629;
	#10 counter$count = 95630;
	#10 counter$count = 95631;
	#10 counter$count = 95632;
	#10 counter$count = 95633;
	#10 counter$count = 95634;
	#10 counter$count = 95635;
	#10 counter$count = 95636;
	#10 counter$count = 95637;
	#10 counter$count = 95638;
	#10 counter$count = 95639;
	#10 counter$count = 95640;
	#10 counter$count = 95641;
	#10 counter$count = 95642;
	#10 counter$count = 95643;
	#10 counter$count = 95644;
	#10 counter$count = 95645;
	#10 counter$count = 95646;
	#10 counter$count = 95647;
	#10 counter$count = 95648;
	#10 counter$count = 95649;
	#10 counter$count = 95650;
	#10 counter$count = 95651;
	#10 counter$count = 95652;
	#10 counter$count = 95653;
	#10 counter$count = 95654;
	#10 counter$count = 95655;
	#10 counter$count = 95656;
	#10 counter$count = 95657;
	#10 counter$count = 95658;
	#10 counter$count = 95659;
	#10 counter$count = 95660;
	#10 counter$count = 95661;
	#10 counter$count = 95662;
	#10 counter$count = 95663;
	#10 counter$count = 95664;
	#10 counter$count = 95665;
	#10 counter$count = 95666;
	#10 counter$count = 95667;
	#10 counter$count = 95668;
	#10 counter$count = 95669;
	#10 counter$count = 95670;
	#10 counter$count = 95671;
	#10 counter$count = 95672;
	#10 counter$count = 95673;
	#10 counter$count = 95674;
	#10 counter$count = 95675;
	#10 counter$count = 95676;
	#10 counter$count = 95677;
	#10 counter$count = 95678;
	#10 counter$count = 95679;
	#10 counter$count = 95680;
	#10 counter$count = 95681;
	#10 counter$count = 95682;
	#10 counter$count = 95683;
	#10 counter$count = 95684;
	#10 counter$count = 95685;
	#10 counter$count = 95686;
	#10 counter$count = 95687;
	#10 counter$count = 95688;
	#10 counter$count = 95689;
	#10 counter$count = 95690;
	#10 counter$count = 95691;
	#10 counter$count = 95692;
	#10 counter$count = 95693;
	#10 counter$count = 95694;
	#10 counter$count = 95695;
	#10 counter$count = 95696;
	#10 counter$count = 95697;
	#10 counter$count = 95698;
	#10 counter$count = 95699;
	#10 counter$count = 95700;
	#10 counter$count = 95701;
	#10 counter$count = 95702;
	#10 counter$count = 95703;
	#10 counter$count = 95704;
	#10 counter$count = 95705;
	#10 counter$count = 95706;
	#10 counter$count = 95707;
	#10 counter$count = 95708;
	#10 counter$count = 95709;
	#10 counter$count = 95710;
	#10 counter$count = 95711;
	#10 counter$count = 95712;
	#10 counter$count = 95713;
	#10 counter$count = 95714;
	#10 counter$count = 95715;
	#10 counter$count = 95716;
	#10 counter$count = 95717;
	#10 counter$count = 95718;
	#10 counter$count = 95719;
	#10 counter$count = 95720;
	#10 counter$count = 95721;
	#10 counter$count = 95722;
	#10 counter$count = 95723;
	#10 counter$count = 95724;
	#10 counter$count = 95725;
	#10 counter$count = 95726;
	#10 counter$count = 95727;
	#10 counter$count = 95728;
	#10 counter$count = 95729;
	#10 counter$count = 95730;
	#10 counter$count = 95731;
	#10 counter$count = 95732;
	#10 counter$count = 95733;
	#10 counter$count = 95734;
	#10 counter$count = 95735;
	#10 counter$count = 95736;
	#10 counter$count = 95737;
	#10 counter$count = 95738;
	#10 counter$count = 95739;
	#10 counter$count = 95740;
	#10 counter$count = 95741;
	#10 counter$count = 95742;
	#10 counter$count = 95743;
	#10 counter$count = 95744;
	#10 counter$count = 95745;
	#10 counter$count = 95746;
	#10 counter$count = 95747;
	#10 counter$count = 95748;
	#10 counter$count = 95749;
	#10 counter$count = 95750;
	#10 counter$count = 95751;
	#10 counter$count = 95752;
	#10 counter$count = 95753;
	#10 counter$count = 95754;
	#10 counter$count = 95755;
	#10 counter$count = 95756;
	#10 counter$count = 95757;
	#10 counter$count = 95758;
	#10 counter$count = 95759;
	#10 counter$count = 95760;
	#10 counter$count = 95761;
	#10 counter$count = 95762;
	#10 counter$count = 95763;
	#10 counter$count = 95764;
	#10 counter$count = 95765;
	#10 counter$count = 95766;
	#10 counter$count = 95767;
	#10 counter$count = 95768;
	#10 counter$count = 95769;
	#10 counter$count = 95770;
	#10 counter$count = 95771;
	#10 counter$count = 95772;
	#10 counter$count = 95773;
	#10 counter$count = 95774;
	#10 counter$count = 95775;
	#10 counter$count = 95776;
	#10 counter$count = 95777;
	#10 counter$count = 95778;
	#10 counter$count = 95779;
	#10 counter$count = 95780;
	#10 counter$count = 95781;
	#10 counter$count = 95782;
	#10 counter$count = 95783;
	#10 counter$count = 95784;
	#10 counter$count = 95785;
	#10 counter$count = 95786;
	#10 counter$count = 95787;
	#10 counter$count = 95788;
	#10 counter$count = 95789;
	#10 counter$count = 95790;
	#10 counter$count = 95791;
	#10 counter$count = 95792;
	#10 counter$count = 95793;
	#10 counter$count = 95794;
	#10 counter$count = 95795;
	#10 counter$count = 95796;
	#10 counter$count = 95797;
	#10 counter$count = 95798;
	#10 counter$count = 95799;
	#10 counter$count = 95800;
	#10 counter$count = 95801;
	#10 counter$count = 95802;
	#10 counter$count = 95803;
	#10 counter$count = 95804;
	#10 counter$count = 95805;
	#10 counter$count = 95806;
	#10 counter$count = 95807;
	#10 counter$count = 95808;
	#10 counter$count = 95809;
	#10 counter$count = 95810;
	#10 counter$count = 95811;
	#10 counter$count = 95812;
	#10 counter$count = 95813;
	#10 counter$count = 95814;
	#10 counter$count = 95815;
	#10 counter$count = 95816;
	#10 counter$count = 95817;
	#10 counter$count = 95818;
	#10 counter$count = 95819;
	#10 counter$count = 95820;
	#10 counter$count = 95821;
	#10 counter$count = 95822;
	#10 counter$count = 95823;
	#10 counter$count = 95824;
	#10 counter$count = 95825;
	#10 counter$count = 95826;
	#10 counter$count = 95827;
	#10 counter$count = 95828;
	#10 counter$count = 95829;
	#10 counter$count = 95830;
	#10 counter$count = 95831;
	#10 counter$count = 95832;
	#10 counter$count = 95833;
	#10 counter$count = 95834;
	#10 counter$count = 95835;
	#10 counter$count = 95836;
	#10 counter$count = 95837;
	#10 counter$count = 95838;
	#10 counter$count = 95839;
	#10 counter$count = 95840;
	#10 counter$count = 95841;
	#10 counter$count = 95842;
	#10 counter$count = 95843;
	#10 counter$count = 95844;
	#10 counter$count = 95845;
	#10 counter$count = 95846;
	#10 counter$count = 95847;
	#10 counter$count = 95848;
	#10 counter$count = 95849;
	#10 counter$count = 95850;
	#10 counter$count = 95851;
	#10 counter$count = 95852;
	#10 counter$count = 95853;
	#10 counter$count = 95854;
	#10 counter$count = 95855;
	#10 counter$count = 95856;
	#10 counter$count = 95857;
	#10 counter$count = 95858;
	#10 counter$count = 95859;
	#10 counter$count = 95860;
	#10 counter$count = 95861;
	#10 counter$count = 95862;
	#10 counter$count = 95863;
	#10 counter$count = 95864;
	#10 counter$count = 95865;
	#10 counter$count = 95866;
	#10 counter$count = 95867;
	#10 counter$count = 95868;
	#10 counter$count = 95869;
	#10 counter$count = 95870;
	#10 counter$count = 95871;
	#10 counter$count = 95872;
	#10 counter$count = 95873;
	#10 counter$count = 95874;
	#10 counter$count = 95875;
	#10 counter$count = 95876;
	#10 counter$count = 95877;
	#10 counter$count = 95878;
	#10 counter$count = 95879;
	#10 counter$count = 95880;
	#10 counter$count = 95881;
	#10 counter$count = 95882;
	#10 counter$count = 95883;
	#10 counter$count = 95884;
	#10 counter$count = 95885;
	#10 counter$count = 95886;
	#10 counter$count = 95887;
	#10 counter$count = 95888;
	#10 counter$count = 95889;
	#10 counter$count = 95890;
	#10 counter$count = 95891;
	#10 counter$count = 95892;
	#10 counter$count = 95893;
	#10 counter$count = 95894;
	#10 counter$count = 95895;
	#10 counter$count = 95896;
	#10 counter$count = 95897;
	#10 counter$count = 95898;
	#10 counter$count = 95899;
	#10 counter$count = 95900;
	#10 counter$count = 95901;
	#10 counter$count = 95902;
	#10 counter$count = 95903;
	#10 counter$count = 95904;
	#10 counter$count = 95905;
	#10 counter$count = 95906;
	#10 counter$count = 95907;
	#10 counter$count = 95908;
	#10 counter$count = 95909;
	#10 counter$count = 95910;
	#10 counter$count = 95911;
	#10 counter$count = 95912;
	#10 counter$count = 95913;
	#10 counter$count = 95914;
	#10 counter$count = 95915;
	#10 counter$count = 95916;
	#10 counter$count = 95917;
	#10 counter$count = 95918;
	#10 counter$count = 95919;
	#10 counter$count = 95920;
	#10 counter$count = 95921;
	#10 counter$count = 95922;
	#10 counter$count = 95923;
	#10 counter$count = 95924;
	#10 counter$count = 95925;
	#10 counter$count = 95926;
	#10 counter$count = 95927;
	#10 counter$count = 95928;
	#10 counter$count = 95929;
	#10 counter$count = 95930;
	#10 counter$count = 95931;
	#10 counter$count = 95932;
	#10 counter$count = 95933;
	#10 counter$count = 95934;
	#10 counter$count = 95935;
	#10 counter$count = 95936;
	#10 counter$count = 95937;
	#10 counter$count = 95938;
	#10 counter$count = 95939;
	#10 counter$count = 95940;
	#10 counter$count = 95941;
	#10 counter$count = 95942;
	#10 counter$count = 95943;
	#10 counter$count = 95944;
	#10 counter$count = 95945;
	#10 counter$count = 95946;
	#10 counter$count = 95947;
	#10 counter$count = 95948;
	#10 counter$count = 95949;
	#10 counter$count = 95950;
	#10 counter$count = 95951;
	#10 counter$count = 95952;
	#10 counter$count = 95953;
	#10 counter$count = 95954;
	#10 counter$count = 95955;
	#10 counter$count = 95956;
	#10 counter$count = 95957;
	#10 counter$count = 95958;
	#10 counter$count = 95959;
	#10 counter$count = 95960;
	#10 counter$count = 95961;
	#10 counter$count = 95962;
	#10 counter$count = 95963;
	#10 counter$count = 95964;
	#10 counter$count = 95965;
	#10 counter$count = 95966;
	#10 counter$count = 95967;
	#10 counter$count = 95968;
	#10 counter$count = 95969;
	#10 counter$count = 95970;
	#10 counter$count = 95971;
	#10 counter$count = 95972;
	#10 counter$count = 95973;
	#10 counter$count = 95974;
	#10 counter$count = 95975;
	#10 counter$count = 95976;
	#10 counter$count = 95977;
	#10 counter$count = 95978;
	#10 counter$count = 95979;
	#10 counter$count = 95980;
	#10 counter$count = 95981;
	#10 counter$count = 95982;
	#10 counter$count = 95983;
	#10 counter$count = 95984;
	#10 counter$count = 95985;
	#10 counter$count = 95986;
	#10 counter$count = 95987;
	#10 counter$count = 95988;
	#10 counter$count = 95989;
	#10 counter$count = 95990;
	#10 counter$count = 95991;
	#10 counter$count = 95992;
	#10 counter$count = 95993;
	#10 counter$count = 95994;
	#10 counter$count = 95995;
	#10 counter$count = 95996;
	#10 counter$count = 95997;
	#10 counter$count = 95998;
	#10 counter$count = 95999;
	#10 counter$count = 96000;
	#10 counter$count = 96001;
	#10 counter$count = 96002;
	#10 counter$count = 96003;
	#10 counter$count = 96004;
	#10 counter$count = 96005;
	#10 counter$count = 96006;
	#10 counter$count = 96007;
	#10 counter$count = 96008;
	#10 counter$count = 96009;
	#10 counter$count = 96010;
	#10 counter$count = 96011;
	#10 counter$count = 96012;
	#10 counter$count = 96013;
	#10 counter$count = 96014;
	#10 counter$count = 96015;
	#10 counter$count = 96016;
	#10 counter$count = 96017;
	#10 counter$count = 96018;
	#10 counter$count = 96019;
	#10 counter$count = 96020;
	#10 counter$count = 96021;
	#10 counter$count = 96022;
	#10 counter$count = 96023;
	#10 counter$count = 96024;
	#10 counter$count = 96025;
	#10 counter$count = 96026;
	#10 counter$count = 96027;
	#10 counter$count = 96028;
	#10 counter$count = 96029;
	#10 counter$count = 96030;
	#10 counter$count = 96031;
	#10 counter$count = 96032;
	#10 counter$count = 96033;
	#10 counter$count = 96034;
	#10 counter$count = 96035;
	#10 counter$count = 96036;
	#10 counter$count = 96037;
	#10 counter$count = 96038;
	#10 counter$count = 96039;
	#10 counter$count = 96040;
	#10 counter$count = 96041;
	#10 counter$count = 96042;
	#10 counter$count = 96043;
	#10 counter$count = 96044;
	#10 counter$count = 96045;
	#10 counter$count = 96046;
	#10 counter$count = 96047;
	#10 counter$count = 96048;
	#10 counter$count = 96049;
	#10 counter$count = 96050;
	#10 counter$count = 96051;
	#10 counter$count = 96052;
	#10 counter$count = 96053;
	#10 counter$count = 96054;
	#10 counter$count = 96055;
	#10 counter$count = 96056;
	#10 counter$count = 96057;
	#10 counter$count = 96058;
	#10 counter$count = 96059;
	#10 counter$count = 96060;
	#10 counter$count = 96061;
	#10 counter$count = 96062;
	#10 counter$count = 96063;
	#10 counter$count = 96064;
	#10 counter$count = 96065;
	#10 counter$count = 96066;
	#10 counter$count = 96067;
	#10 counter$count = 96068;
	#10 counter$count = 96069;
	#10 counter$count = 96070;
	#10 counter$count = 96071;
	#10 counter$count = 96072;
	#10 counter$count = 96073;
	#10 counter$count = 96074;
	#10 counter$count = 96075;
	#10 counter$count = 96076;
	#10 counter$count = 96077;
	#10 counter$count = 96078;
	#10 counter$count = 96079;
	#10 counter$count = 96080;
	#10 counter$count = 96081;
	#10 counter$count = 96082;
	#10 counter$count = 96083;
	#10 counter$count = 96084;
	#10 counter$count = 96085;
	#10 counter$count = 96086;
	#10 counter$count = 96087;
	#10 counter$count = 96088;
	#10 counter$count = 96089;
	#10 counter$count = 96090;
	#10 counter$count = 96091;
	#10 counter$count = 96092;
	#10 counter$count = 96093;
	#10 counter$count = 96094;
	#10 counter$count = 96095;
	#10 counter$count = 96096;
	#10 counter$count = 96097;
	#10 counter$count = 96098;
	#10 counter$count = 96099;
	#10 counter$count = 96100;
	#10 counter$count = 96101;
	#10 counter$count = 96102;
	#10 counter$count = 96103;
	#10 counter$count = 96104;
	#10 counter$count = 96105;
	#10 counter$count = 96106;
	#10 counter$count = 96107;
	#10 counter$count = 96108;
	#10 counter$count = 96109;
	#10 counter$count = 96110;
	#10 counter$count = 96111;
	#10 counter$count = 96112;
	#10 counter$count = 96113;
	#10 counter$count = 96114;
	#10 counter$count = 96115;
	#10 counter$count = 96116;
	#10 counter$count = 96117;
	#10 counter$count = 96118;
	#10 counter$count = 96119;
	#10 counter$count = 96120;
	#10 counter$count = 96121;
	#10 counter$count = 96122;
	#10 counter$count = 96123;
	#10 counter$count = 96124;
	#10 counter$count = 96125;
	#10 counter$count = 96126;
	#10 counter$count = 96127;
	#10 counter$count = 96128;
	#10 counter$count = 96129;
	#10 counter$count = 96130;
	#10 counter$count = 96131;
	#10 counter$count = 96132;
	#10 counter$count = 96133;
	#10 counter$count = 96134;
	#10 counter$count = 96135;
	#10 counter$count = 96136;
	#10 counter$count = 96137;
	#10 counter$count = 96138;
	#10 counter$count = 96139;
	#10 counter$count = 96140;
	#10 counter$count = 96141;
	#10 counter$count = 96142;
	#10 counter$count = 96143;
	#10 counter$count = 96144;
	#10 counter$count = 96145;
	#10 counter$count = 96146;
	#10 counter$count = 96147;
	#10 counter$count = 96148;
	#10 counter$count = 96149;
	#10 counter$count = 96150;
	#10 counter$count = 96151;
	#10 counter$count = 96152;
	#10 counter$count = 96153;
	#10 counter$count = 96154;
	#10 counter$count = 96155;
	#10 counter$count = 96156;
	#10 counter$count = 96157;
	#10 counter$count = 96158;
	#10 counter$count = 96159;
	#10 counter$count = 96160;
	#10 counter$count = 96161;
	#10 counter$count = 96162;
	#10 counter$count = 96163;
	#10 counter$count = 96164;
	#10 counter$count = 96165;
	#10 counter$count = 96166;
	#10 counter$count = 96167;
	#10 counter$count = 96168;
	#10 counter$count = 96169;
	#10 counter$count = 96170;
	#10 counter$count = 96171;
	#10 counter$count = 96172;
	#10 counter$count = 96173;
	#10 counter$count = 96174;
	#10 counter$count = 96175;
	#10 counter$count = 96176;
	#10 counter$count = 96177;
	#10 counter$count = 96178;
	#10 counter$count = 96179;
	#10 counter$count = 96180;
	#10 counter$count = 96181;
	#10 counter$count = 96182;
	#10 counter$count = 96183;
	#10 counter$count = 96184;
	#10 counter$count = 96185;
	#10 counter$count = 96186;
	#10 counter$count = 96187;
	#10 counter$count = 96188;
	#10 counter$count = 96189;
	#10 counter$count = 96190;
	#10 counter$count = 96191;
	#10 counter$count = 96192;
	#10 counter$count = 96193;
	#10 counter$count = 96194;
	#10 counter$count = 96195;
	#10 counter$count = 96196;
	#10 counter$count = 96197;
	#10 counter$count = 96198;
	#10 counter$count = 96199;
	#10 counter$count = 96200;
	#10 counter$count = 96201;
	#10 counter$count = 96202;
	#10 counter$count = 96203;
	#10 counter$count = 96204;
	#10 counter$count = 96205;
	#10 counter$count = 96206;
	#10 counter$count = 96207;
	#10 counter$count = 96208;
	#10 counter$count = 96209;
	#10 counter$count = 96210;
	#10 counter$count = 96211;
	#10 counter$count = 96212;
	#10 counter$count = 96213;
	#10 counter$count = 96214;
	#10 counter$count = 96215;
	#10 counter$count = 96216;
	#10 counter$count = 96217;
	#10 counter$count = 96218;
	#10 counter$count = 96219;
	#10 counter$count = 96220;
	#10 counter$count = 96221;
	#10 counter$count = 96222;
	#10 counter$count = 96223;
	#10 counter$count = 96224;
	#10 counter$count = 96225;
	#10 counter$count = 96226;
	#10 counter$count = 96227;
	#10 counter$count = 96228;
	#10 counter$count = 96229;
	#10 counter$count = 96230;
	#10 counter$count = 96231;
	#10 counter$count = 96232;
	#10 counter$count = 96233;
	#10 counter$count = 96234;
	#10 counter$count = 96235;
	#10 counter$count = 96236;
	#10 counter$count = 96237;
	#10 counter$count = 96238;
	#10 counter$count = 96239;
	#10 counter$count = 96240;
	#10 counter$count = 96241;
	#10 counter$count = 96242;
	#10 counter$count = 96243;
	#10 counter$count = 96244;
	#10 counter$count = 96245;
	#10 counter$count = 96246;
	#10 counter$count = 96247;
	#10 counter$count = 96248;
	#10 counter$count = 96249;
	#10 counter$count = 96250;
	#10 counter$count = 96251;
	#10 counter$count = 96252;
	#10 counter$count = 96253;
	#10 counter$count = 96254;
	#10 counter$count = 96255;
	#10 counter$count = 96256;
	#10 counter$count = 96257;
	#10 counter$count = 96258;
	#10 counter$count = 96259;
	#10 counter$count = 96260;
	#10 counter$count = 96261;
	#10 counter$count = 96262;
	#10 counter$count = 96263;
	#10 counter$count = 96264;
	#10 counter$count = 96265;
	#10 counter$count = 96266;
	#10 counter$count = 96267;
	#10 counter$count = 96268;
	#10 counter$count = 96269;
	#10 counter$count = 96270;
	#10 counter$count = 96271;
	#10 counter$count = 96272;
	#10 counter$count = 96273;
	#10 counter$count = 96274;
	#10 counter$count = 96275;
	#10 counter$count = 96276;
	#10 counter$count = 96277;
	#10 counter$count = 96278;
	#10 counter$count = 96279;
	#10 counter$count = 96280;
	#10 counter$count = 96281;
	#10 counter$count = 96282;
	#10 counter$count = 96283;
	#10 counter$count = 96284;
	#10 counter$count = 96285;
	#10 counter$count = 96286;
	#10 counter$count = 96287;
	#10 counter$count = 96288;
	#10 counter$count = 96289;
	#10 counter$count = 96290;
	#10 counter$count = 96291;
	#10 counter$count = 96292;
	#10 counter$count = 96293;
	#10 counter$count = 96294;
	#10 counter$count = 96295;
	#10 counter$count = 96296;
	#10 counter$count = 96297;
	#10 counter$count = 96298;
	#10 counter$count = 96299;
	#10 counter$count = 96300;
	#10 counter$count = 96301;
	#10 counter$count = 96302;
	#10 counter$count = 96303;
	#10 counter$count = 96304;
	#10 counter$count = 96305;
	#10 counter$count = 96306;
	#10 counter$count = 96307;
	#10 counter$count = 96308;
	#10 counter$count = 96309;
	#10 counter$count = 96310;
	#10 counter$count = 96311;
	#10 counter$count = 96312;
	#10 counter$count = 96313;
	#10 counter$count = 96314;
	#10 counter$count = 96315;
	#10 counter$count = 96316;
	#10 counter$count = 96317;
	#10 counter$count = 96318;
	#10 counter$count = 96319;
	#10 counter$count = 96320;
	#10 counter$count = 96321;
	#10 counter$count = 96322;
	#10 counter$count = 96323;
	#10 counter$count = 96324;
	#10 counter$count = 96325;
	#10 counter$count = 96326;
	#10 counter$count = 96327;
	#10 counter$count = 96328;
	#10 counter$count = 96329;
	#10 counter$count = 96330;
	#10 counter$count = 96331;
	#10 counter$count = 96332;
	#10 counter$count = 96333;
	#10 counter$count = 96334;
	#10 counter$count = 96335;
	#10 counter$count = 96336;
	#10 counter$count = 96337;
	#10 counter$count = 96338;
	#10 counter$count = 96339;
	#10 counter$count = 96340;
	#10 counter$count = 96341;
	#10 counter$count = 96342;
	#10 counter$count = 96343;
	#10 counter$count = 96344;
	#10 counter$count = 96345;
	#10 counter$count = 96346;
	#10 counter$count = 96347;
	#10 counter$count = 96348;
	#10 counter$count = 96349;
	#10 counter$count = 96350;
	#10 counter$count = 96351;
	#10 counter$count = 96352;
	#10 counter$count = 96353;
	#10 counter$count = 96354;
	#10 counter$count = 96355;
	#10 counter$count = 96356;
	#10 counter$count = 96357;
	#10 counter$count = 96358;
	#10 counter$count = 96359;
	#10 counter$count = 96360;
	#10 counter$count = 96361;
	#10 counter$count = 96362;
	#10 counter$count = 96363;
	#10 counter$count = 96364;
	#10 counter$count = 96365;
	#10 counter$count = 96366;
	#10 counter$count = 96367;
	#10 counter$count = 96368;
	#10 counter$count = 96369;
	#10 counter$count = 96370;
	#10 counter$count = 96371;
	#10 counter$count = 96372;
	#10 counter$count = 96373;
	#10 counter$count = 96374;
	#10 counter$count = 96375;
	#10 counter$count = 96376;
	#10 counter$count = 96377;
	#10 counter$count = 96378;
	#10 counter$count = 96379;
	#10 counter$count = 96380;
	#10 counter$count = 96381;
	#10 counter$count = 96382;
	#10 counter$count = 96383;
	#10 counter$count = 96384;
	#10 counter$count = 96385;
	#10 counter$count = 96386;
	#10 counter$count = 96387;
	#10 counter$count = 96388;
	#10 counter$count = 96389;
	#10 counter$count = 96390;
	#10 counter$count = 96391;
	#10 counter$count = 96392;
	#10 counter$count = 96393;
	#10 counter$count = 96394;
	#10 counter$count = 96395;
	#10 counter$count = 96396;
	#10 counter$count = 96397;
	#10 counter$count = 96398;
	#10 counter$count = 96399;
	#10 counter$count = 96400;
	#10 counter$count = 96401;
	#10 counter$count = 96402;
	#10 counter$count = 96403;
	#10 counter$count = 96404;
	#10 counter$count = 96405;
	#10 counter$count = 96406;
	#10 counter$count = 96407;
	#10 counter$count = 96408;
	#10 counter$count = 96409;
	#10 counter$count = 96410;
	#10 counter$count = 96411;
	#10 counter$count = 96412;
	#10 counter$count = 96413;
	#10 counter$count = 96414;
	#10 counter$count = 96415;
	#10 counter$count = 96416;
	#10 counter$count = 96417;
	#10 counter$count = 96418;
	#10 counter$count = 96419;
	#10 counter$count = 96420;
	#10 counter$count = 96421;
	#10 counter$count = 96422;
	#10 counter$count = 96423;
	#10 counter$count = 96424;
	#10 counter$count = 96425;
	#10 counter$count = 96426;
	#10 counter$count = 96427;
	#10 counter$count = 96428;
	#10 counter$count = 96429;
	#10 counter$count = 96430;
	#10 counter$count = 96431;
	#10 counter$count = 96432;
	#10 counter$count = 96433;
	#10 counter$count = 96434;
	#10 counter$count = 96435;
	#10 counter$count = 96436;
	#10 counter$count = 96437;
	#10 counter$count = 96438;
	#10 counter$count = 96439;
	#10 counter$count = 96440;
	#10 counter$count = 96441;
	#10 counter$count = 96442;
	#10 counter$count = 96443;
	#10 counter$count = 96444;
	#10 counter$count = 96445;
	#10 counter$count = 96446;
	#10 counter$count = 96447;
	#10 counter$count = 96448;
	#10 counter$count = 96449;
	#10 counter$count = 96450;
	#10 counter$count = 96451;
	#10 counter$count = 96452;
	#10 counter$count = 96453;
	#10 counter$count = 96454;
	#10 counter$count = 96455;
	#10 counter$count = 96456;
	#10 counter$count = 96457;
	#10 counter$count = 96458;
	#10 counter$count = 96459;
	#10 counter$count = 96460;
	#10 counter$count = 96461;
	#10 counter$count = 96462;
	#10 counter$count = 96463;
	#10 counter$count = 96464;
	#10 counter$count = 96465;
	#10 counter$count = 96466;
	#10 counter$count = 96467;
	#10 counter$count = 96468;
	#10 counter$count = 96469;
	#10 counter$count = 96470;
	#10 counter$count = 96471;
	#10 counter$count = 96472;
	#10 counter$count = 96473;
	#10 counter$count = 96474;
	#10 counter$count = 96475;
	#10 counter$count = 96476;
	#10 counter$count = 96477;
	#10 counter$count = 96478;
	#10 counter$count = 96479;
	#10 counter$count = 96480;
	#10 counter$count = 96481;
	#10 counter$count = 96482;
	#10 counter$count = 96483;
	#10 counter$count = 96484;
	#10 counter$count = 96485;
	#10 counter$count = 96486;
	#10 counter$count = 96487;
	#10 counter$count = 96488;
	#10 counter$count = 96489;
	#10 counter$count = 96490;
	#10 counter$count = 96491;
	#10 counter$count = 96492;
	#10 counter$count = 96493;
	#10 counter$count = 96494;
	#10 counter$count = 96495;
	#10 counter$count = 96496;
	#10 counter$count = 96497;
	#10 counter$count = 96498;
	#10 counter$count = 96499;
	#10 counter$count = 96500;
	#10 counter$count = 96501;
	#10 counter$count = 96502;
	#10 counter$count = 96503;
	#10 counter$count = 96504;
	#10 counter$count = 96505;
	#10 counter$count = 96506;
	#10 counter$count = 96507;
	#10 counter$count = 96508;
	#10 counter$count = 96509;
	#10 counter$count = 96510;
	#10 counter$count = 96511;
	#10 counter$count = 96512;
	#10 counter$count = 96513;
	#10 counter$count = 96514;
	#10 counter$count = 96515;
	#10 counter$count = 96516;
	#10 counter$count = 96517;
	#10 counter$count = 96518;
	#10 counter$count = 96519;
	#10 counter$count = 96520;
	#10 counter$count = 96521;
	#10 counter$count = 96522;
	#10 counter$count = 96523;
	#10 counter$count = 96524;
	#10 counter$count = 96525;
	#10 counter$count = 96526;
	#10 counter$count = 96527;
	#10 counter$count = 96528;
	#10 counter$count = 96529;
	#10 counter$count = 96530;
	#10 counter$count = 96531;
	#10 counter$count = 96532;
	#10 counter$count = 96533;
	#10 counter$count = 96534;
	#10 counter$count = 96535;
	#10 counter$count = 96536;
	#10 counter$count = 96537;
	#10 counter$count = 96538;
	#10 counter$count = 96539;
	#10 counter$count = 96540;
	#10 counter$count = 96541;
	#10 counter$count = 96542;
	#10 counter$count = 96543;
	#10 counter$count = 96544;
	#10 counter$count = 96545;
	#10 counter$count = 96546;
	#10 counter$count = 96547;
	#10 counter$count = 96548;
	#10 counter$count = 96549;
	#10 counter$count = 96550;
	#10 counter$count = 96551;
	#10 counter$count = 96552;
	#10 counter$count = 96553;
	#10 counter$count = 96554;
	#10 counter$count = 96555;
	#10 counter$count = 96556;
	#10 counter$count = 96557;
	#10 counter$count = 96558;
	#10 counter$count = 96559;
	#10 counter$count = 96560;
	#10 counter$count = 96561;
	#10 counter$count = 96562;
	#10 counter$count = 96563;
	#10 counter$count = 96564;
	#10 counter$count = 96565;
	#10 counter$count = 96566;
	#10 counter$count = 96567;
	#10 counter$count = 96568;
	#10 counter$count = 96569;
	#10 counter$count = 96570;
	#10 counter$count = 96571;
	#10 counter$count = 96572;
	#10 counter$count = 96573;
	#10 counter$count = 96574;
	#10 counter$count = 96575;
	#10 counter$count = 96576;
	#10 counter$count = 96577;
	#10 counter$count = 96578;
	#10 counter$count = 96579;
	#10 counter$count = 96580;
	#10 counter$count = 96581;
	#10 counter$count = 96582;
	#10 counter$count = 96583;
	#10 counter$count = 96584;
	#10 counter$count = 96585;
	#10 counter$count = 96586;
	#10 counter$count = 96587;
	#10 counter$count = 96588;
	#10 counter$count = 96589;
	#10 counter$count = 96590;
	#10 counter$count = 96591;
	#10 counter$count = 96592;
	#10 counter$count = 96593;
	#10 counter$count = 96594;
	#10 counter$count = 96595;
	#10 counter$count = 96596;
	#10 counter$count = 96597;
	#10 counter$count = 96598;
	#10 counter$count = 96599;
	#10 counter$count = 96600;
	#10 counter$count = 96601;
	#10 counter$count = 96602;
	#10 counter$count = 96603;
	#10 counter$count = 96604;
	#10 counter$count = 96605;
	#10 counter$count = 96606;
	#10 counter$count = 96607;
	#10 counter$count = 96608;
	#10 counter$count = 96609;
	#10 counter$count = 96610;
	#10 counter$count = 96611;
	#10 counter$count = 96612;
	#10 counter$count = 96613;
	#10 counter$count = 96614;
	#10 counter$count = 96615;
	#10 counter$count = 96616;
	#10 counter$count = 96617;
	#10 counter$count = 96618;
	#10 counter$count = 96619;
	#10 counter$count = 96620;
	#10 counter$count = 96621;
	#10 counter$count = 96622;
	#10 counter$count = 96623;
	#10 counter$count = 96624;
	#10 counter$count = 96625;
	#10 counter$count = 96626;
	#10 counter$count = 96627;
	#10 counter$count = 96628;
	#10 counter$count = 96629;
	#10 counter$count = 96630;
	#10 counter$count = 96631;
	#10 counter$count = 96632;
	#10 counter$count = 96633;
	#10 counter$count = 96634;
	#10 counter$count = 96635;
	#10 counter$count = 96636;
	#10 counter$count = 96637;
	#10 counter$count = 96638;
	#10 counter$count = 96639;
	#10 counter$count = 96640;
	#10 counter$count = 96641;
	#10 counter$count = 96642;
	#10 counter$count = 96643;
	#10 counter$count = 96644;
	#10 counter$count = 96645;
	#10 counter$count = 96646;
	#10 counter$count = 96647;
	#10 counter$count = 96648;
	#10 counter$count = 96649;
	#10 counter$count = 96650;
	#10 counter$count = 96651;
	#10 counter$count = 96652;
	#10 counter$count = 96653;
	#10 counter$count = 96654;
	#10 counter$count = 96655;
	#10 counter$count = 96656;
	#10 counter$count = 96657;
	#10 counter$count = 96658;
	#10 counter$count = 96659;
	#10 counter$count = 96660;
	#10 counter$count = 96661;
	#10 counter$count = 96662;
	#10 counter$count = 96663;
	#10 counter$count = 96664;
	#10 counter$count = 96665;
	#10 counter$count = 96666;
	#10 counter$count = 96667;
	#10 counter$count = 96668;
	#10 counter$count = 96669;
	#10 counter$count = 96670;
	#10 counter$count = 96671;
	#10 counter$count = 96672;
	#10 counter$count = 96673;
	#10 counter$count = 96674;
	#10 counter$count = 96675;
	#10 counter$count = 96676;
	#10 counter$count = 96677;
	#10 counter$count = 96678;
	#10 counter$count = 96679;
	#10 counter$count = 96680;
	#10 counter$count = 96681;
	#10 counter$count = 96682;
	#10 counter$count = 96683;
	#10 counter$count = 96684;
	#10 counter$count = 96685;
	#10 counter$count = 96686;
	#10 counter$count = 96687;
	#10 counter$count = 96688;
	#10 counter$count = 96689;
	#10 counter$count = 96690;
	#10 counter$count = 96691;
	#10 counter$count = 96692;
	#10 counter$count = 96693;
	#10 counter$count = 96694;
	#10 counter$count = 96695;
	#10 counter$count = 96696;
	#10 counter$count = 96697;
	#10 counter$count = 96698;
	#10 counter$count = 96699;
	#10 counter$count = 96700;
	#10 counter$count = 96701;
	#10 counter$count = 96702;
	#10 counter$count = 96703;
	#10 counter$count = 96704;
	#10 counter$count = 96705;
	#10 counter$count = 96706;
	#10 counter$count = 96707;
	#10 counter$count = 96708;
	#10 counter$count = 96709;
	#10 counter$count = 96710;
	#10 counter$count = 96711;
	#10 counter$count = 96712;
	#10 counter$count = 96713;
	#10 counter$count = 96714;
	#10 counter$count = 96715;
	#10 counter$count = 96716;
	#10 counter$count = 96717;
	#10 counter$count = 96718;
	#10 counter$count = 96719;
	#10 counter$count = 96720;
	#10 counter$count = 96721;
	#10 counter$count = 96722;
	#10 counter$count = 96723;
	#10 counter$count = 96724;
	#10 counter$count = 96725;
	#10 counter$count = 96726;
	#10 counter$count = 96727;
	#10 counter$count = 96728;
	#10 counter$count = 96729;
	#10 counter$count = 96730;
	#10 counter$count = 96731;
	#10 counter$count = 96732;
	#10 counter$count = 96733;
	#10 counter$count = 96734;
	#10 counter$count = 96735;
	#10 counter$count = 96736;
	#10 counter$count = 96737;
	#10 counter$count = 96738;
	#10 counter$count = 96739;
	#10 counter$count = 96740;
	#10 counter$count = 96741;
	#10 counter$count = 96742;
	#10 counter$count = 96743;
	#10 counter$count = 96744;
	#10 counter$count = 96745;
	#10 counter$count = 96746;
	#10 counter$count = 96747;
	#10 counter$count = 96748;
	#10 counter$count = 96749;
	#10 counter$count = 96750;
	#10 counter$count = 96751;
	#10 counter$count = 96752;
	#10 counter$count = 96753;
	#10 counter$count = 96754;
	#10 counter$count = 96755;
	#10 counter$count = 96756;
	#10 counter$count = 96757;
	#10 counter$count = 96758;
	#10 counter$count = 96759;
	#10 counter$count = 96760;
	#10 counter$count = 96761;
	#10 counter$count = 96762;
	#10 counter$count = 96763;
	#10 counter$count = 96764;
	#10 counter$count = 96765;
	#10 counter$count = 96766;
	#10 counter$count = 96767;
	#10 counter$count = 96768;
	#10 counter$count = 96769;
	#10 counter$count = 96770;
	#10 counter$count = 96771;
	#10 counter$count = 96772;
	#10 counter$count = 96773;
	#10 counter$count = 96774;
	#10 counter$count = 96775;
	#10 counter$count = 96776;
	#10 counter$count = 96777;
	#10 counter$count = 96778;
	#10 counter$count = 96779;
	#10 counter$count = 96780;
	#10 counter$count = 96781;
	#10 counter$count = 96782;
	#10 counter$count = 96783;
	#10 counter$count = 96784;
	#10 counter$count = 96785;
	#10 counter$count = 96786;
	#10 counter$count = 96787;
	#10 counter$count = 96788;
	#10 counter$count = 96789;
	#10 counter$count = 96790;
	#10 counter$count = 96791;
	#10 counter$count = 96792;
	#10 counter$count = 96793;
	#10 counter$count = 96794;
	#10 counter$count = 96795;
	#10 counter$count = 96796;
	#10 counter$count = 96797;
	#10 counter$count = 96798;
	#10 counter$count = 96799;
	#10 counter$count = 96800;
	#10 counter$count = 96801;
	#10 counter$count = 96802;
	#10 counter$count = 96803;
	#10 counter$count = 96804;
	#10 counter$count = 96805;
	#10 counter$count = 96806;
	#10 counter$count = 96807;
	#10 counter$count = 96808;
	#10 counter$count = 96809;
	#10 counter$count = 96810;
	#10 counter$count = 96811;
	#10 counter$count = 96812;
	#10 counter$count = 96813;
	#10 counter$count = 96814;
	#10 counter$count = 96815;
	#10 counter$count = 96816;
	#10 counter$count = 96817;
	#10 counter$count = 96818;
	#10 counter$count = 96819;
	#10 counter$count = 96820;
	#10 counter$count = 96821;
	#10 counter$count = 96822;
	#10 counter$count = 96823;
	#10 counter$count = 96824;
	#10 counter$count = 96825;
	#10 counter$count = 96826;
	#10 counter$count = 96827;
	#10 counter$count = 96828;
	#10 counter$count = 96829;
	#10 counter$count = 96830;
	#10 counter$count = 96831;
	#10 counter$count = 96832;
	#10 counter$count = 96833;
	#10 counter$count = 96834;
	#10 counter$count = 96835;
	#10 counter$count = 96836;
	#10 counter$count = 96837;
	#10 counter$count = 96838;
	#10 counter$count = 96839;
	#10 counter$count = 96840;
	#10 counter$count = 96841;
	#10 counter$count = 96842;
	#10 counter$count = 96843;
	#10 counter$count = 96844;
	#10 counter$count = 96845;
	#10 counter$count = 96846;
	#10 counter$count = 96847;
	#10 counter$count = 96848;
	#10 counter$count = 96849;
	#10 counter$count = 96850;
	#10 counter$count = 96851;
	#10 counter$count = 96852;
	#10 counter$count = 96853;
	#10 counter$count = 96854;
	#10 counter$count = 96855;
	#10 counter$count = 96856;
	#10 counter$count = 96857;
	#10 counter$count = 96858;
	#10 counter$count = 96859;
	#10 counter$count = 96860;
	#10 counter$count = 96861;
	#10 counter$count = 96862;
	#10 counter$count = 96863;
	#10 counter$count = 96864;
	#10 counter$count = 96865;
	#10 counter$count = 96866;
	#10 counter$count = 96867;
	#10 counter$count = 96868;
	#10 counter$count = 96869;
	#10 counter$count = 96870;
	#10 counter$count = 96871;
	#10 counter$count = 96872;
	#10 counter$count = 96873;
	#10 counter$count = 96874;
	#10 counter$count = 96875;
	#10 counter$count = 96876;
	#10 counter$count = 96877;
	#10 counter$count = 96878;
	#10 counter$count = 96879;
	#10 counter$count = 96880;
	#10 counter$count = 96881;
	#10 counter$count = 96882;
	#10 counter$count = 96883;
	#10 counter$count = 96884;
	#10 counter$count = 96885;
	#10 counter$count = 96886;
	#10 counter$count = 96887;
	#10 counter$count = 96888;
	#10 counter$count = 96889;
	#10 counter$count = 96890;
	#10 counter$count = 96891;
	#10 counter$count = 96892;
	#10 counter$count = 96893;
	#10 counter$count = 96894;
	#10 counter$count = 96895;
	#10 counter$count = 96896;
	#10 counter$count = 96897;
	#10 counter$count = 96898;
	#10 counter$count = 96899;
	#10 counter$count = 96900;
	#10 counter$count = 96901;
	#10 counter$count = 96902;
	#10 counter$count = 96903;
	#10 counter$count = 96904;
	#10 counter$count = 96905;
	#10 counter$count = 96906;
	#10 counter$count = 96907;
	#10 counter$count = 96908;
	#10 counter$count = 96909;
	#10 counter$count = 96910;
	#10 counter$count = 96911;
	#10 counter$count = 96912;
	#10 counter$count = 96913;
	#10 counter$count = 96914;
	#10 counter$count = 96915;
	#10 counter$count = 96916;
	#10 counter$count = 96917;
	#10 counter$count = 96918;
	#10 counter$count = 96919;
	#10 counter$count = 96920;
	#10 counter$count = 96921;
	#10 counter$count = 96922;
	#10 counter$count = 96923;
	#10 counter$count = 96924;
	#10 counter$count = 96925;
	#10 counter$count = 96926;
	#10 counter$count = 96927;
	#10 counter$count = 96928;
	#10 counter$count = 96929;
	#10 counter$count = 96930;
	#10 counter$count = 96931;
	#10 counter$count = 96932;
	#10 counter$count = 96933;
	#10 counter$count = 96934;
	#10 counter$count = 96935;
	#10 counter$count = 96936;
	#10 counter$count = 96937;
	#10 counter$count = 96938;
	#10 counter$count = 96939;
	#10 counter$count = 96940;
	#10 counter$count = 96941;
	#10 counter$count = 96942;
	#10 counter$count = 96943;
	#10 counter$count = 96944;
	#10 counter$count = 96945;
	#10 counter$count = 96946;
	#10 counter$count = 96947;
	#10 counter$count = 96948;
	#10 counter$count = 96949;
	#10 counter$count = 96950;
	#10 counter$count = 96951;
	#10 counter$count = 96952;
	#10 counter$count = 96953;
	#10 counter$count = 96954;
	#10 counter$count = 96955;
	#10 counter$count = 96956;
	#10 counter$count = 96957;
	#10 counter$count = 96958;
	#10 counter$count = 96959;
	#10 counter$count = 96960;
	#10 counter$count = 96961;
	#10 counter$count = 96962;
	#10 counter$count = 96963;
	#10 counter$count = 96964;
	#10 counter$count = 96965;
	#10 counter$count = 96966;
	#10 counter$count = 96967;
	#10 counter$count = 96968;
	#10 counter$count = 96969;
	#10 counter$count = 96970;
	#10 counter$count = 96971;
	#10 counter$count = 96972;
	#10 counter$count = 96973;
	#10 counter$count = 96974;
	#10 counter$count = 96975;
	#10 counter$count = 96976;
	#10 counter$count = 96977;
	#10 counter$count = 96978;
	#10 counter$count = 96979;
	#10 counter$count = 96980;
	#10 counter$count = 96981;
	#10 counter$count = 96982;
	#10 counter$count = 96983;
	#10 counter$count = 96984;
	#10 counter$count = 96985;
	#10 counter$count = 96986;
	#10 counter$count = 96987;
	#10 counter$count = 96988;
	#10 counter$count = 96989;
	#10 counter$count = 96990;
	#10 counter$count = 96991;
	#10 counter$count = 96992;
	#10 counter$count = 96993;
	#10 counter$count = 96994;
	#10 counter$count = 96995;
	#10 counter$count = 96996;
	#10 counter$count = 96997;
	#10 counter$count = 96998;
	#10 counter$count = 96999;
	#10 counter$count = 97000;
	#10 counter$count = 97001;
	#10 counter$count = 97002;
	#10 counter$count = 97003;
	#10 counter$count = 97004;
	#10 counter$count = 97005;
	#10 counter$count = 97006;
	#10 counter$count = 97007;
	#10 counter$count = 97008;
	#10 counter$count = 97009;
	#10 counter$count = 97010;
	#10 counter$count = 97011;
	#10 counter$count = 97012;
	#10 counter$count = 97013;
	#10 counter$count = 97014;
	#10 counter$count = 97015;
	#10 counter$count = 97016;
	#10 counter$count = 97017;
	#10 counter$count = 97018;
	#10 counter$count = 97019;
	#10 counter$count = 97020;
	#10 counter$count = 97021;
	#10 counter$count = 97022;
	#10 counter$count = 97023;
	#10 counter$count = 97024;
	#10 counter$count = 97025;
	#10 counter$count = 97026;
	#10 counter$count = 97027;
	#10 counter$count = 97028;
	#10 counter$count = 97029;
	#10 counter$count = 97030;
	#10 counter$count = 97031;
	#10 counter$count = 97032;
	#10 counter$count = 97033;
	#10 counter$count = 97034;
	#10 counter$count = 97035;
	#10 counter$count = 97036;
	#10 counter$count = 97037;
	#10 counter$count = 97038;
	#10 counter$count = 97039;
	#10 counter$count = 97040;
	#10 counter$count = 97041;
	#10 counter$count = 97042;
	#10 counter$count = 97043;
	#10 counter$count = 97044;
	#10 counter$count = 97045;
	#10 counter$count = 97046;
	#10 counter$count = 97047;
	#10 counter$count = 97048;
	#10 counter$count = 97049;
	#10 counter$count = 97050;
	#10 counter$count = 97051;
	#10 counter$count = 97052;
	#10 counter$count = 97053;
	#10 counter$count = 97054;
	#10 counter$count = 97055;
	#10 counter$count = 97056;
	#10 counter$count = 97057;
	#10 counter$count = 97058;
	#10 counter$count = 97059;
	#10 counter$count = 97060;
	#10 counter$count = 97061;
	#10 counter$count = 97062;
	#10 counter$count = 97063;
	#10 counter$count = 97064;
	#10 counter$count = 97065;
	#10 counter$count = 97066;
	#10 counter$count = 97067;
	#10 counter$count = 97068;
	#10 counter$count = 97069;
	#10 counter$count = 97070;
	#10 counter$count = 97071;
	#10 counter$count = 97072;
	#10 counter$count = 97073;
	#10 counter$count = 97074;
	#10 counter$count = 97075;
	#10 counter$count = 97076;
	#10 counter$count = 97077;
	#10 counter$count = 97078;
	#10 counter$count = 97079;
	#10 counter$count = 97080;
	#10 counter$count = 97081;
	#10 counter$count = 97082;
	#10 counter$count = 97083;
	#10 counter$count = 97084;
	#10 counter$count = 97085;
	#10 counter$count = 97086;
	#10 counter$count = 97087;
	#10 counter$count = 97088;
	#10 counter$count = 97089;
	#10 counter$count = 97090;
	#10 counter$count = 97091;
	#10 counter$count = 97092;
	#10 counter$count = 97093;
	#10 counter$count = 97094;
	#10 counter$count = 97095;
	#10 counter$count = 97096;
	#10 counter$count = 97097;
	#10 counter$count = 97098;
	#10 counter$count = 97099;
	#10 counter$count = 97100;
	#10 counter$count = 97101;
	#10 counter$count = 97102;
	#10 counter$count = 97103;
	#10 counter$count = 97104;
	#10 counter$count = 97105;
	#10 counter$count = 97106;
	#10 counter$count = 97107;
	#10 counter$count = 97108;
	#10 counter$count = 97109;
	#10 counter$count = 97110;
	#10 counter$count = 97111;
	#10 counter$count = 97112;
	#10 counter$count = 97113;
	#10 counter$count = 97114;
	#10 counter$count = 97115;
	#10 counter$count = 97116;
	#10 counter$count = 97117;
	#10 counter$count = 97118;
	#10 counter$count = 97119;
	#10 counter$count = 97120;
	#10 counter$count = 97121;
	#10 counter$count = 97122;
	#10 counter$count = 97123;
	#10 counter$count = 97124;
	#10 counter$count = 97125;
	#10 counter$count = 97126;
	#10 counter$count = 97127;
	#10 counter$count = 97128;
	#10 counter$count = 97129;
	#10 counter$count = 97130;
	#10 counter$count = 97131;
	#10 counter$count = 97132;
	#10 counter$count = 97133;
	#10 counter$count = 97134;
	#10 counter$count = 97135;
	#10 counter$count = 97136;
	#10 counter$count = 97137;
	#10 counter$count = 97138;
	#10 counter$count = 97139;
	#10 counter$count = 97140;
	#10 counter$count = 97141;
	#10 counter$count = 97142;
	#10 counter$count = 97143;
	#10 counter$count = 97144;
	#10 counter$count = 97145;
	#10 counter$count = 97146;
	#10 counter$count = 97147;
	#10 counter$count = 97148;
	#10 counter$count = 97149;
	#10 counter$count = 97150;
	#10 counter$count = 97151;
	#10 counter$count = 97152;
	#10 counter$count = 97153;
	#10 counter$count = 97154;
	#10 counter$count = 97155;
	#10 counter$count = 97156;
	#10 counter$count = 97157;
	#10 counter$count = 97158;
	#10 counter$count = 97159;
	#10 counter$count = 97160;
	#10 counter$count = 97161;
	#10 counter$count = 97162;
	#10 counter$count = 97163;
	#10 counter$count = 97164;
	#10 counter$count = 97165;
	#10 counter$count = 97166;
	#10 counter$count = 97167;
	#10 counter$count = 97168;
	#10 counter$count = 97169;
	#10 counter$count = 97170;
	#10 counter$count = 97171;
	#10 counter$count = 97172;
	#10 counter$count = 97173;
	#10 counter$count = 97174;
	#10 counter$count = 97175;
	#10 counter$count = 97176;
	#10 counter$count = 97177;
	#10 counter$count = 97178;
	#10 counter$count = 97179;
	#10 counter$count = 97180;
	#10 counter$count = 97181;
	#10 counter$count = 97182;
	#10 counter$count = 97183;
	#10 counter$count = 97184;
	#10 counter$count = 97185;
	#10 counter$count = 97186;
	#10 counter$count = 97187;
	#10 counter$count = 97188;
	#10 counter$count = 97189;
	#10 counter$count = 97190;
	#10 counter$count = 97191;
	#10 counter$count = 97192;
	#10 counter$count = 97193;
	#10 counter$count = 97194;
	#10 counter$count = 97195;
	#10 counter$count = 97196;
	#10 counter$count = 97197;
	#10 counter$count = 97198;
	#10 counter$count = 97199;
	#10 counter$count = 97200;
	#10 counter$count = 97201;
	#10 counter$count = 97202;
	#10 counter$count = 97203;
	#10 counter$count = 97204;
	#10 counter$count = 97205;
	#10 counter$count = 97206;
	#10 counter$count = 97207;
	#10 counter$count = 97208;
	#10 counter$count = 97209;
	#10 counter$count = 97210;
	#10 counter$count = 97211;
	#10 counter$count = 97212;
	#10 counter$count = 97213;
	#10 counter$count = 97214;
	#10 counter$count = 97215;
	#10 counter$count = 97216;
	#10 counter$count = 97217;
	#10 counter$count = 97218;
	#10 counter$count = 97219;
	#10 counter$count = 97220;
	#10 counter$count = 97221;
	#10 counter$count = 97222;
	#10 counter$count = 97223;
	#10 counter$count = 97224;
	#10 counter$count = 97225;
	#10 counter$count = 97226;
	#10 counter$count = 97227;
	#10 counter$count = 97228;
	#10 counter$count = 97229;
	#10 counter$count = 97230;
	#10 counter$count = 97231;
	#10 counter$count = 97232;
	#10 counter$count = 97233;
	#10 counter$count = 97234;
	#10 counter$count = 97235;
	#10 counter$count = 97236;
	#10 counter$count = 97237;
	#10 counter$count = 97238;
	#10 counter$count = 97239;
	#10 counter$count = 97240;
	#10 counter$count = 97241;
	#10 counter$count = 97242;
	#10 counter$count = 97243;
	#10 counter$count = 97244;
	#10 counter$count = 97245;
	#10 counter$count = 97246;
	#10 counter$count = 97247;
	#10 counter$count = 97248;
	#10 counter$count = 97249;
	#10 counter$count = 97250;
	#10 counter$count = 97251;
	#10 counter$count = 97252;
	#10 counter$count = 97253;
	#10 counter$count = 97254;
	#10 counter$count = 97255;
	#10 counter$count = 97256;
	#10 counter$count = 97257;
	#10 counter$count = 97258;
	#10 counter$count = 97259;
	#10 counter$count = 97260;
	#10 counter$count = 97261;
	#10 counter$count = 97262;
	#10 counter$count = 97263;
	#10 counter$count = 97264;
	#10 counter$count = 97265;
	#10 counter$count = 97266;
	#10 counter$count = 97267;
	#10 counter$count = 97268;
	#10 counter$count = 97269;
	#10 counter$count = 97270;
	#10 counter$count = 97271;
	#10 counter$count = 97272;
	#10 counter$count = 97273;
	#10 counter$count = 97274;
	#10 counter$count = 97275;
	#10 counter$count = 97276;
	#10 counter$count = 97277;
	#10 counter$count = 97278;
	#10 counter$count = 97279;
	#10 counter$count = 97280;
	#10 counter$count = 97281;
	#10 counter$count = 97282;
	#10 counter$count = 97283;
	#10 counter$count = 97284;
	#10 counter$count = 97285;
	#10 counter$count = 97286;
	#10 counter$count = 97287;
	#10 counter$count = 97288;
	#10 counter$count = 97289;
	#10 counter$count = 97290;
	#10 counter$count = 97291;
	#10 counter$count = 97292;
	#10 counter$count = 97293;
	#10 counter$count = 97294;
	#10 counter$count = 97295;
	#10 counter$count = 97296;
	#10 counter$count = 97297;
	#10 counter$count = 97298;
	#10 counter$count = 97299;
	#10 counter$count = 97300;
	#10 counter$count = 97301;
	#10 counter$count = 97302;
	#10 counter$count = 97303;
	#10 counter$count = 97304;
	#10 counter$count = 97305;
	#10 counter$count = 97306;
	#10 counter$count = 97307;
	#10 counter$count = 97308;
	#10 counter$count = 97309;
	#10 counter$count = 97310;
	#10 counter$count = 97311;
	#10 counter$count = 97312;
	#10 counter$count = 97313;
	#10 counter$count = 97314;
	#10 counter$count = 97315;
	#10 counter$count = 97316;
	#10 counter$count = 97317;
	#10 counter$count = 97318;
	#10 counter$count = 97319;
	#10 counter$count = 97320;
	#10 counter$count = 97321;
	#10 counter$count = 97322;
	#10 counter$count = 97323;
	#10 counter$count = 97324;
	#10 counter$count = 97325;
	#10 counter$count = 97326;
	#10 counter$count = 97327;
	#10 counter$count = 97328;
	#10 counter$count = 97329;
	#10 counter$count = 97330;
	#10 counter$count = 97331;
	#10 counter$count = 97332;
	#10 counter$count = 97333;
	#10 counter$count = 97334;
	#10 counter$count = 97335;
	#10 counter$count = 97336;
	#10 counter$count = 97337;
	#10 counter$count = 97338;
	#10 counter$count = 97339;
	#10 counter$count = 97340;
	#10 counter$count = 97341;
	#10 counter$count = 97342;
	#10 counter$count = 97343;
	#10 counter$count = 97344;
	#10 counter$count = 97345;
	#10 counter$count = 97346;
	#10 counter$count = 97347;
	#10 counter$count = 97348;
	#10 counter$count = 97349;
	#10 counter$count = 97350;
	#10 counter$count = 97351;
	#10 counter$count = 97352;
	#10 counter$count = 97353;
	#10 counter$count = 97354;
	#10 counter$count = 97355;
	#10 counter$count = 97356;
	#10 counter$count = 97357;
	#10 counter$count = 97358;
	#10 counter$count = 97359;
	#10 counter$count = 97360;
	#10 counter$count = 97361;
	#10 counter$count = 97362;
	#10 counter$count = 97363;
	#10 counter$count = 97364;
	#10 counter$count = 97365;
	#10 counter$count = 97366;
	#10 counter$count = 97367;
	#10 counter$count = 97368;
	#10 counter$count = 97369;
	#10 counter$count = 97370;
	#10 counter$count = 97371;
	#10 counter$count = 97372;
	#10 counter$count = 97373;
	#10 counter$count = 97374;
	#10 counter$count = 97375;
	#10 counter$count = 97376;
	#10 counter$count = 97377;
	#10 counter$count = 97378;
	#10 counter$count = 97379;
	#10 counter$count = 97380;
	#10 counter$count = 97381;
	#10 counter$count = 97382;
	#10 counter$count = 97383;
	#10 counter$count = 97384;
	#10 counter$count = 97385;
	#10 counter$count = 97386;
	#10 counter$count = 97387;
	#10 counter$count = 97388;
	#10 counter$count = 97389;
	#10 counter$count = 97390;
	#10 counter$count = 97391;
	#10 counter$count = 97392;
	#10 counter$count = 97393;
	#10 counter$count = 97394;
	#10 counter$count = 97395;
	#10 counter$count = 97396;
	#10 counter$count = 97397;
	#10 counter$count = 97398;
	#10 counter$count = 97399;
	#10 counter$count = 97400;
	#10 counter$count = 97401;
	#10 counter$count = 97402;
	#10 counter$count = 97403;
	#10 counter$count = 97404;
	#10 counter$count = 97405;
	#10 counter$count = 97406;
	#10 counter$count = 97407;
	#10 counter$count = 97408;
	#10 counter$count = 97409;
	#10 counter$count = 97410;
	#10 counter$count = 97411;
	#10 counter$count = 97412;
	#10 counter$count = 97413;
	#10 counter$count = 97414;
	#10 counter$count = 97415;
	#10 counter$count = 97416;
	#10 counter$count = 97417;
	#10 counter$count = 97418;
	#10 counter$count = 97419;
	#10 counter$count = 97420;
	#10 counter$count = 97421;
	#10 counter$count = 97422;
	#10 counter$count = 97423;
	#10 counter$count = 97424;
	#10 counter$count = 97425;
	#10 counter$count = 97426;
	#10 counter$count = 97427;
	#10 counter$count = 97428;
	#10 counter$count = 97429;
	#10 counter$count = 97430;
	#10 counter$count = 97431;
	#10 counter$count = 97432;
	#10 counter$count = 97433;
	#10 counter$count = 97434;
	#10 counter$count = 97435;
	#10 counter$count = 97436;
	#10 counter$count = 97437;
	#10 counter$count = 97438;
	#10 counter$count = 97439;
	#10 counter$count = 97440;
	#10 counter$count = 97441;
	#10 counter$count = 97442;
	#10 counter$count = 97443;
	#10 counter$count = 97444;
	#10 counter$count = 97445;
	#10 counter$count = 97446;
	#10 counter$count = 97447;
	#10 counter$count = 97448;
	#10 counter$count = 97449;
	#10 counter$count = 97450;
	#10 counter$count = 97451;
	#10 counter$count = 97452;
	#10 counter$count = 97453;
	#10 counter$count = 97454;
	#10 counter$count = 97455;
	#10 counter$count = 97456;
	#10 counter$count = 97457;
	#10 counter$count = 97458;
	#10 counter$count = 97459;
	#10 counter$count = 97460;
	#10 counter$count = 97461;
	#10 counter$count = 97462;
	#10 counter$count = 97463;
	#10 counter$count = 97464;
	#10 counter$count = 97465;
	#10 counter$count = 97466;
	#10 counter$count = 97467;
	#10 counter$count = 97468;
	#10 counter$count = 97469;
	#10 counter$count = 97470;
	#10 counter$count = 97471;
	#10 counter$count = 97472;
	#10 counter$count = 97473;
	#10 counter$count = 97474;
	#10 counter$count = 97475;
	#10 counter$count = 97476;
	#10 counter$count = 97477;
	#10 counter$count = 97478;
	#10 counter$count = 97479;
	#10 counter$count = 97480;
	#10 counter$count = 97481;
	#10 counter$count = 97482;
	#10 counter$count = 97483;
	#10 counter$count = 97484;
	#10 counter$count = 97485;
	#10 counter$count = 97486;
	#10 counter$count = 97487;
	#10 counter$count = 97488;
	#10 counter$count = 97489;
	#10 counter$count = 97490;
	#10 counter$count = 97491;
	#10 counter$count = 97492;
	#10 counter$count = 97493;
	#10 counter$count = 97494;
	#10 counter$count = 97495;
	#10 counter$count = 97496;
	#10 counter$count = 97497;
	#10 counter$count = 97498;
	#10 counter$count = 97499;
	#10 counter$count = 97500;
	#10 counter$count = 97501;
	#10 counter$count = 97502;
	#10 counter$count = 97503;
	#10 counter$count = 97504;
	#10 counter$count = 97505;
	#10 counter$count = 97506;
	#10 counter$count = 97507;
	#10 counter$count = 97508;
	#10 counter$count = 97509;
	#10 counter$count = 97510;
	#10 counter$count = 97511;
	#10 counter$count = 97512;
	#10 counter$count = 97513;
	#10 counter$count = 97514;
	#10 counter$count = 97515;
	#10 counter$count = 97516;
	#10 counter$count = 97517;
	#10 counter$count = 97518;
	#10 counter$count = 97519;
	#10 counter$count = 97520;
	#10 counter$count = 97521;
	#10 counter$count = 97522;
	#10 counter$count = 97523;
	#10 counter$count = 97524;
	#10 counter$count = 97525;
	#10 counter$count = 97526;
	#10 counter$count = 97527;
	#10 counter$count = 97528;
	#10 counter$count = 97529;
	#10 counter$count = 97530;
	#10 counter$count = 97531;
	#10 counter$count = 97532;
	#10 counter$count = 97533;
	#10 counter$count = 97534;
	#10 counter$count = 97535;
	#10 counter$count = 97536;
	#10 counter$count = 97537;
	#10 counter$count = 97538;
	#10 counter$count = 97539;
	#10 counter$count = 97540;
	#10 counter$count = 97541;
	#10 counter$count = 97542;
	#10 counter$count = 97543;
	#10 counter$count = 97544;
	#10 counter$count = 97545;
	#10 counter$count = 97546;
	#10 counter$count = 97547;
	#10 counter$count = 97548;
	#10 counter$count = 97549;
	#10 counter$count = 97550;
	#10 counter$count = 97551;
	#10 counter$count = 97552;
	#10 counter$count = 97553;
	#10 counter$count = 97554;
	#10 counter$count = 97555;
	#10 counter$count = 97556;
	#10 counter$count = 97557;
	#10 counter$count = 97558;
	#10 counter$count = 97559;
	#10 counter$count = 97560;
	#10 counter$count = 97561;
	#10 counter$count = 97562;
	#10 counter$count = 97563;
	#10 counter$count = 97564;
	#10 counter$count = 97565;
	#10 counter$count = 97566;
	#10 counter$count = 97567;
	#10 counter$count = 97568;
	#10 counter$count = 97569;
	#10 counter$count = 97570;
	#10 counter$count = 97571;
	#10 counter$count = 97572;
	#10 counter$count = 97573;
	#10 counter$count = 97574;
	#10 counter$count = 97575;
	#10 counter$count = 97576;
	#10 counter$count = 97577;
	#10 counter$count = 97578;
	#10 counter$count = 97579;
	#10 counter$count = 97580;
	#10 counter$count = 97581;
	#10 counter$count = 97582;
	#10 counter$count = 97583;
	#10 counter$count = 97584;
	#10 counter$count = 97585;
	#10 counter$count = 97586;
	#10 counter$count = 97587;
	#10 counter$count = 97588;
	#10 counter$count = 97589;
	#10 counter$count = 97590;
	#10 counter$count = 97591;
	#10 counter$count = 97592;
	#10 counter$count = 97593;
	#10 counter$count = 97594;
	#10 counter$count = 97595;
	#10 counter$count = 97596;
	#10 counter$count = 97597;
	#10 counter$count = 97598;
	#10 counter$count = 97599;
	#10 counter$count = 97600;
	#10 counter$count = 97601;
	#10 counter$count = 97602;
	#10 counter$count = 97603;
	#10 counter$count = 97604;
	#10 counter$count = 97605;
	#10 counter$count = 97606;
	#10 counter$count = 97607;
	#10 counter$count = 97608;
	#10 counter$count = 97609;
	#10 counter$count = 97610;
	#10 counter$count = 97611;
	#10 counter$count = 97612;
	#10 counter$count = 97613;
	#10 counter$count = 97614;
	#10 counter$count = 97615;
	#10 counter$count = 97616;
	#10 counter$count = 97617;
	#10 counter$count = 97618;
	#10 counter$count = 97619;
	#10 counter$count = 97620;
	#10 counter$count = 97621;
	#10 counter$count = 97622;
	#10 counter$count = 97623;
	#10 counter$count = 97624;
	#10 counter$count = 97625;
	#10 counter$count = 97626;
	#10 counter$count = 97627;
	#10 counter$count = 97628;
	#10 counter$count = 97629;
	#10 counter$count = 97630;
	#10 counter$count = 97631;
	#10 counter$count = 97632;
	#10 counter$count = 97633;
	#10 counter$count = 97634;
	#10 counter$count = 97635;
	#10 counter$count = 97636;
	#10 counter$count = 97637;
	#10 counter$count = 97638;
	#10 counter$count = 97639;
	#10 counter$count = 97640;
	#10 counter$count = 97641;
	#10 counter$count = 97642;
	#10 counter$count = 97643;
	#10 counter$count = 97644;
	#10 counter$count = 97645;
	#10 counter$count = 97646;
	#10 counter$count = 97647;
	#10 counter$count = 97648;
	#10 counter$count = 97649;
	#10 counter$count = 97650;
	#10 counter$count = 97651;
	#10 counter$count = 97652;
	#10 counter$count = 97653;
	#10 counter$count = 97654;
	#10 counter$count = 97655;
	#10 counter$count = 97656;
	#10 counter$count = 97657;
	#10 counter$count = 97658;
	#10 counter$count = 97659;
	#10 counter$count = 97660;
	#10 counter$count = 97661;
	#10 counter$count = 97662;
	#10 counter$count = 97663;
	#10 counter$count = 97664;
	#10 counter$count = 97665;
	#10 counter$count = 97666;
	#10 counter$count = 97667;
	#10 counter$count = 97668;
	#10 counter$count = 97669;
	#10 counter$count = 97670;
	#10 counter$count = 97671;
	#10 counter$count = 97672;
	#10 counter$count = 97673;
	#10 counter$count = 97674;
	#10 counter$count = 97675;
	#10 counter$count = 97676;
	#10 counter$count = 97677;
	#10 counter$count = 97678;
	#10 counter$count = 97679;
	#10 counter$count = 97680;
	#10 counter$count = 97681;
	#10 counter$count = 97682;
	#10 counter$count = 97683;
	#10 counter$count = 97684;
	#10 counter$count = 97685;
	#10 counter$count = 97686;
	#10 counter$count = 97687;
	#10 counter$count = 97688;
	#10 counter$count = 97689;
	#10 counter$count = 97690;
	#10 counter$count = 97691;
	#10 counter$count = 97692;
	#10 counter$count = 97693;
	#10 counter$count = 97694;
	#10 counter$count = 97695;
	#10 counter$count = 97696;
	#10 counter$count = 97697;
	#10 counter$count = 97698;
	#10 counter$count = 97699;
	#10 counter$count = 97700;
	#10 counter$count = 97701;
	#10 counter$count = 97702;
	#10 counter$count = 97703;
	#10 counter$count = 97704;
	#10 counter$count = 97705;
	#10 counter$count = 97706;
	#10 counter$count = 97707;
	#10 counter$count = 97708;
	#10 counter$count = 97709;
	#10 counter$count = 97710;
	#10 counter$count = 97711;
	#10 counter$count = 97712;
	#10 counter$count = 97713;
	#10 counter$count = 97714;
	#10 counter$count = 97715;
	#10 counter$count = 97716;
	#10 counter$count = 97717;
	#10 counter$count = 97718;
	#10 counter$count = 97719;
	#10 counter$count = 97720;
	#10 counter$count = 97721;
	#10 counter$count = 97722;
	#10 counter$count = 97723;
	#10 counter$count = 97724;
	#10 counter$count = 97725;
	#10 counter$count = 97726;
	#10 counter$count = 97727;
	#10 counter$count = 97728;
	#10 counter$count = 97729;
	#10 counter$count = 97730;
	#10 counter$count = 97731;
	#10 counter$count = 97732;
	#10 counter$count = 97733;
	#10 counter$count = 97734;
	#10 counter$count = 97735;
	#10 counter$count = 97736;
	#10 counter$count = 97737;
	#10 counter$count = 97738;
	#10 counter$count = 97739;
	#10 counter$count = 97740;
	#10 counter$count = 97741;
	#10 counter$count = 97742;
	#10 counter$count = 97743;
	#10 counter$count = 97744;
	#10 counter$count = 97745;
	#10 counter$count = 97746;
	#10 counter$count = 97747;
	#10 counter$count = 97748;
	#10 counter$count = 97749;
	#10 counter$count = 97750;
	#10 counter$count = 97751;
	#10 counter$count = 97752;
	#10 counter$count = 97753;
	#10 counter$count = 97754;
	#10 counter$count = 97755;
	#10 counter$count = 97756;
	#10 counter$count = 97757;
	#10 counter$count = 97758;
	#10 counter$count = 97759;
	#10 counter$count = 97760;
	#10 counter$count = 97761;
	#10 counter$count = 97762;
	#10 counter$count = 97763;
	#10 counter$count = 97764;
	#10 counter$count = 97765;
	#10 counter$count = 97766;
	#10 counter$count = 97767;
	#10 counter$count = 97768;
	#10 counter$count = 97769;
	#10 counter$count = 97770;
	#10 counter$count = 97771;
	#10 counter$count = 97772;
	#10 counter$count = 97773;
	#10 counter$count = 97774;
	#10 counter$count = 97775;
	#10 counter$count = 97776;
	#10 counter$count = 97777;
	#10 counter$count = 97778;
	#10 counter$count = 97779;
	#10 counter$count = 97780;
	#10 counter$count = 97781;
	#10 counter$count = 97782;
	#10 counter$count = 97783;
	#10 counter$count = 97784;
	#10 counter$count = 97785;
	#10 counter$count = 97786;
	#10 counter$count = 97787;
	#10 counter$count = 97788;
	#10 counter$count = 97789;
	#10 counter$count = 97790;
	#10 counter$count = 97791;
	#10 counter$count = 97792;
	#10 counter$count = 97793;
	#10 counter$count = 97794;
	#10 counter$count = 97795;
	#10 counter$count = 97796;
	#10 counter$count = 97797;
	#10 counter$count = 97798;
	#10 counter$count = 97799;
	#10 counter$count = 97800;
	#10 counter$count = 97801;
	#10 counter$count = 97802;
	#10 counter$count = 97803;
	#10 counter$count = 97804;
	#10 counter$count = 97805;
	#10 counter$count = 97806;
	#10 counter$count = 97807;
	#10 counter$count = 97808;
	#10 counter$count = 97809;
	#10 counter$count = 97810;
	#10 counter$count = 97811;
	#10 counter$count = 97812;
	#10 counter$count = 97813;
	#10 counter$count = 97814;
	#10 counter$count = 97815;
	#10 counter$count = 97816;
	#10 counter$count = 97817;
	#10 counter$count = 97818;
	#10 counter$count = 97819;
	#10 counter$count = 97820;
	#10 counter$count = 97821;
	#10 counter$count = 97822;
	#10 counter$count = 97823;
	#10 counter$count = 97824;
	#10 counter$count = 97825;
	#10 counter$count = 97826;
	#10 counter$count = 97827;
	#10 counter$count = 97828;
	#10 counter$count = 97829;
	#10 counter$count = 97830;
	#10 counter$count = 97831;
	#10 counter$count = 97832;
	#10 counter$count = 97833;
	#10 counter$count = 97834;
	#10 counter$count = 97835;
	#10 counter$count = 97836;
	#10 counter$count = 97837;
	#10 counter$count = 97838;
	#10 counter$count = 97839;
	#10 counter$count = 97840;
	#10 counter$count = 97841;
	#10 counter$count = 97842;
	#10 counter$count = 97843;
	#10 counter$count = 97844;
	#10 counter$count = 97845;
	#10 counter$count = 97846;
	#10 counter$count = 97847;
	#10 counter$count = 97848;
	#10 counter$count = 97849;
	#10 counter$count = 97850;
	#10 counter$count = 97851;
	#10 counter$count = 97852;
	#10 counter$count = 97853;
	#10 counter$count = 97854;
	#10 counter$count = 97855;
	#10 counter$count = 97856;
	#10 counter$count = 97857;
	#10 counter$count = 97858;
	#10 counter$count = 97859;
	#10 counter$count = 97860;
	#10 counter$count = 97861;
	#10 counter$count = 97862;
	#10 counter$count = 97863;
	#10 counter$count = 97864;
	#10 counter$count = 97865;
	#10 counter$count = 97866;
	#10 counter$count = 97867;
	#10 counter$count = 97868;
	#10 counter$count = 97869;
	#10 counter$count = 97870;
	#10 counter$count = 97871;
	#10 counter$count = 97872;
	#10 counter$count = 97873;
	#10 counter$count = 97874;
	#10 counter$count = 97875;
	#10 counter$count = 97876;
	#10 counter$count = 97877;
	#10 counter$count = 97878;
	#10 counter$count = 97879;
	#10 counter$count = 97880;
	#10 counter$count = 97881;
	#10 counter$count = 97882;
	#10 counter$count = 97883;
	#10 counter$count = 97884;
	#10 counter$count = 97885;
	#10 counter$count = 97886;
	#10 counter$count = 97887;
	#10 counter$count = 97888;
	#10 counter$count = 97889;
	#10 counter$count = 97890;
	#10 counter$count = 97891;
	#10 counter$count = 97892;
	#10 counter$count = 97893;
	#10 counter$count = 97894;
	#10 counter$count = 97895;
	#10 counter$count = 97896;
	#10 counter$count = 97897;
	#10 counter$count = 97898;
	#10 counter$count = 97899;
	#10 counter$count = 97900;
	#10 counter$count = 97901;
	#10 counter$count = 97902;
	#10 counter$count = 97903;
	#10 counter$count = 97904;
	#10 counter$count = 97905;
	#10 counter$count = 97906;
	#10 counter$count = 97907;
	#10 counter$count = 97908;
	#10 counter$count = 97909;
	#10 counter$count = 97910;
	#10 counter$count = 97911;
	#10 counter$count = 97912;
	#10 counter$count = 97913;
	#10 counter$count = 97914;
	#10 counter$count = 97915;
	#10 counter$count = 97916;
	#10 counter$count = 97917;
	#10 counter$count = 97918;
	#10 counter$count = 97919;
	#10 counter$count = 97920;
	#10 counter$count = 97921;
	#10 counter$count = 97922;
	#10 counter$count = 97923;
	#10 counter$count = 97924;
	#10 counter$count = 97925;
	#10 counter$count = 97926;
	#10 counter$count = 97927;
	#10 counter$count = 97928;
	#10 counter$count = 97929;
	#10 counter$count = 97930;
	#10 counter$count = 97931;
	#10 counter$count = 97932;
	#10 counter$count = 97933;
	#10 counter$count = 97934;
	#10 counter$count = 97935;
	#10 counter$count = 97936;
	#10 counter$count = 97937;
	#10 counter$count = 97938;
	#10 counter$count = 97939;
	#10 counter$count = 97940;
	#10 counter$count = 97941;
	#10 counter$count = 97942;
	#10 counter$count = 97943;
	#10 counter$count = 97944;
	#10 counter$count = 97945;
	#10 counter$count = 97946;
	#10 counter$count = 97947;
	#10 counter$count = 97948;
	#10 counter$count = 97949;
	#10 counter$count = 97950;
	#10 counter$count = 97951;
	#10 counter$count = 97952;
	#10 counter$count = 97953;
	#10 counter$count = 97954;
	#10 counter$count = 97955;
	#10 counter$count = 97956;
	#10 counter$count = 97957;
	#10 counter$count = 97958;
	#10 counter$count = 97959;
	#10 counter$count = 97960;
	#10 counter$count = 97961;
	#10 counter$count = 97962;
	#10 counter$count = 97963;
	#10 counter$count = 97964;
	#10 counter$count = 97965;
	#10 counter$count = 97966;
	#10 counter$count = 97967;
	#10 counter$count = 97968;
	#10 counter$count = 97969;
	#10 counter$count = 97970;
	#10 counter$count = 97971;
	#10 counter$count = 97972;
	#10 counter$count = 97973;
	#10 counter$count = 97974;
	#10 counter$count = 97975;
	#10 counter$count = 97976;
	#10 counter$count = 97977;
	#10 counter$count = 97978;
	#10 counter$count = 97979;
	#10 counter$count = 97980;
	#10 counter$count = 97981;
	#10 counter$count = 97982;
	#10 counter$count = 97983;
	#10 counter$count = 97984;
	#10 counter$count = 97985;
	#10 counter$count = 97986;
	#10 counter$count = 97987;
	#10 counter$count = 97988;
	#10 counter$count = 97989;
	#10 counter$count = 97990;
	#10 counter$count = 97991;
	#10 counter$count = 97992;
	#10 counter$count = 97993;
	#10 counter$count = 97994;
	#10 counter$count = 97995;
	#10 counter$count = 97996;
	#10 counter$count = 97997;
	#10 counter$count = 97998;
	#10 counter$count = 97999;
	#10 counter$count = 98000;
	#10 counter$count = 98001;
	#10 counter$count = 98002;
	#10 counter$count = 98003;
	#10 counter$count = 98004;
	#10 counter$count = 98005;
	#10 counter$count = 98006;
	#10 counter$count = 98007;
	#10 counter$count = 98008;
	#10 counter$count = 98009;
	#10 counter$count = 98010;
	#10 counter$count = 98011;
	#10 counter$count = 98012;
	#10 counter$count = 98013;
	#10 counter$count = 98014;
	#10 counter$count = 98015;
	#10 counter$count = 98016;
	#10 counter$count = 98017;
	#10 counter$count = 98018;
	#10 counter$count = 98019;
	#10 counter$count = 98020;
	#10 counter$count = 98021;
	#10 counter$count = 98022;
	#10 counter$count = 98023;
	#10 counter$count = 98024;
	#10 counter$count = 98025;
	#10 counter$count = 98026;
	#10 counter$count = 98027;
	#10 counter$count = 98028;
	#10 counter$count = 98029;
	#10 counter$count = 98030;
	#10 counter$count = 98031;
	#10 counter$count = 98032;
	#10 counter$count = 98033;
	#10 counter$count = 98034;
	#10 counter$count = 98035;
	#10 counter$count = 98036;
	#10 counter$count = 98037;
	#10 counter$count = 98038;
	#10 counter$count = 98039;
	#10 counter$count = 98040;
	#10 counter$count = 98041;
	#10 counter$count = 98042;
	#10 counter$count = 98043;
	#10 counter$count = 98044;
	#10 counter$count = 98045;
	#10 counter$count = 98046;
	#10 counter$count = 98047;
	#10 counter$count = 98048;
	#10 counter$count = 98049;
	#10 counter$count = 98050;
	#10 counter$count = 98051;
	#10 counter$count = 98052;
	#10 counter$count = 98053;
	#10 counter$count = 98054;
	#10 counter$count = 98055;
	#10 counter$count = 98056;
	#10 counter$count = 98057;
	#10 counter$count = 98058;
	#10 counter$count = 98059;
	#10 counter$count = 98060;
	#10 counter$count = 98061;
	#10 counter$count = 98062;
	#10 counter$count = 98063;
	#10 counter$count = 98064;
	#10 counter$count = 98065;
	#10 counter$count = 98066;
	#10 counter$count = 98067;
	#10 counter$count = 98068;
	#10 counter$count = 98069;
	#10 counter$count = 98070;
	#10 counter$count = 98071;
	#10 counter$count = 98072;
	#10 counter$count = 98073;
	#10 counter$count = 98074;
	#10 counter$count = 98075;
	#10 counter$count = 98076;
	#10 counter$count = 98077;
	#10 counter$count = 98078;
	#10 counter$count = 98079;
	#10 counter$count = 98080;
	#10 counter$count = 98081;
	#10 counter$count = 98082;
	#10 counter$count = 98083;
	#10 counter$count = 98084;
	#10 counter$count = 98085;
	#10 counter$count = 98086;
	#10 counter$count = 98087;
	#10 counter$count = 98088;
	#10 counter$count = 98089;
	#10 counter$count = 98090;
	#10 counter$count = 98091;
	#10 counter$count = 98092;
	#10 counter$count = 98093;
	#10 counter$count = 98094;
	#10 counter$count = 98095;
	#10 counter$count = 98096;
	#10 counter$count = 98097;
	#10 counter$count = 98098;
	#10 counter$count = 98099;
	#10 counter$count = 98100;
	#10 counter$count = 98101;
	#10 counter$count = 98102;
	#10 counter$count = 98103;
	#10 counter$count = 98104;
	#10 counter$count = 98105;
	#10 counter$count = 98106;
	#10 counter$count = 98107;
	#10 counter$count = 98108;
	#10 counter$count = 98109;
	#10 counter$count = 98110;
	#10 counter$count = 98111;
	#10 counter$count = 98112;
	#10 counter$count = 98113;
	#10 counter$count = 98114;
	#10 counter$count = 98115;
	#10 counter$count = 98116;
	#10 counter$count = 98117;
	#10 counter$count = 98118;
	#10 counter$count = 98119;
	#10 counter$count = 98120;
	#10 counter$count = 98121;
	#10 counter$count = 98122;
	#10 counter$count = 98123;
	#10 counter$count = 98124;
	#10 counter$count = 98125;
	#10 counter$count = 98126;
	#10 counter$count = 98127;
	#10 counter$count = 98128;
	#10 counter$count = 98129;
	#10 counter$count = 98130;
	#10 counter$count = 98131;
	#10 counter$count = 98132;
	#10 counter$count = 98133;
	#10 counter$count = 98134;
	#10 counter$count = 98135;
	#10 counter$count = 98136;
	#10 counter$count = 98137;
	#10 counter$count = 98138;
	#10 counter$count = 98139;
	#10 counter$count = 98140;
	#10 counter$count = 98141;
	#10 counter$count = 98142;
	#10 counter$count = 98143;
	#10 counter$count = 98144;
	#10 counter$count = 98145;
	#10 counter$count = 98146;
	#10 counter$count = 98147;
	#10 counter$count = 98148;
	#10 counter$count = 98149;
	#10 counter$count = 98150;
	#10 counter$count = 98151;
	#10 counter$count = 98152;
	#10 counter$count = 98153;
	#10 counter$count = 98154;
	#10 counter$count = 98155;
	#10 counter$count = 98156;
	#10 counter$count = 98157;
	#10 counter$count = 98158;
	#10 counter$count = 98159;
	#10 counter$count = 98160;
	#10 counter$count = 98161;
	#10 counter$count = 98162;
	#10 counter$count = 98163;
	#10 counter$count = 98164;
	#10 counter$count = 98165;
	#10 counter$count = 98166;
	#10 counter$count = 98167;
	#10 counter$count = 98168;
	#10 counter$count = 98169;
	#10 counter$count = 98170;
	#10 counter$count = 98171;
	#10 counter$count = 98172;
	#10 counter$count = 98173;
	#10 counter$count = 98174;
	#10 counter$count = 98175;
	#10 counter$count = 98176;
	#10 counter$count = 98177;
	#10 counter$count = 98178;
	#10 counter$count = 98179;
	#10 counter$count = 98180;
	#10 counter$count = 98181;
	#10 counter$count = 98182;
	#10 counter$count = 98183;
	#10 counter$count = 98184;
	#10 counter$count = 98185;
	#10 counter$count = 98186;
	#10 counter$count = 98187;
	#10 counter$count = 98188;
	#10 counter$count = 98189;
	#10 counter$count = 98190;
	#10 counter$count = 98191;
	#10 counter$count = 98192;
	#10 counter$count = 98193;
	#10 counter$count = 98194;
	#10 counter$count = 98195;
	#10 counter$count = 98196;
	#10 counter$count = 98197;
	#10 counter$count = 98198;
	#10 counter$count = 98199;
	#10 counter$count = 98200;
	#10 counter$count = 98201;
	#10 counter$count = 98202;
	#10 counter$count = 98203;
	#10 counter$count = 98204;
	#10 counter$count = 98205;
	#10 counter$count = 98206;
	#10 counter$count = 98207;
	#10 counter$count = 98208;
	#10 counter$count = 98209;
	#10 counter$count = 98210;
	#10 counter$count = 98211;
	#10 counter$count = 98212;
	#10 counter$count = 98213;
	#10 counter$count = 98214;
	#10 counter$count = 98215;
	#10 counter$count = 98216;
	#10 counter$count = 98217;
	#10 counter$count = 98218;
	#10 counter$count = 98219;
	#10 counter$count = 98220;
	#10 counter$count = 98221;
	#10 counter$count = 98222;
	#10 counter$count = 98223;
	#10 counter$count = 98224;
	#10 counter$count = 98225;
	#10 counter$count = 98226;
	#10 counter$count = 98227;
	#10 counter$count = 98228;
	#10 counter$count = 98229;
	#10 counter$count = 98230;
	#10 counter$count = 98231;
	#10 counter$count = 98232;
	#10 counter$count = 98233;
	#10 counter$count = 98234;
	#10 counter$count = 98235;
	#10 counter$count = 98236;
	#10 counter$count = 98237;
	#10 counter$count = 98238;
	#10 counter$count = 98239;
	#10 counter$count = 98240;
	#10 counter$count = 98241;
	#10 counter$count = 98242;
	#10 counter$count = 98243;
	#10 counter$count = 98244;
	#10 counter$count = 98245;
	#10 counter$count = 98246;
	#10 counter$count = 98247;
	#10 counter$count = 98248;
	#10 counter$count = 98249;
	#10 counter$count = 98250;
	#10 counter$count = 98251;
	#10 counter$count = 98252;
	#10 counter$count = 98253;
	#10 counter$count = 98254;
	#10 counter$count = 98255;
	#10 counter$count = 98256;
	#10 counter$count = 98257;
	#10 counter$count = 98258;
	#10 counter$count = 98259;
	#10 counter$count = 98260;
	#10 counter$count = 98261;
	#10 counter$count = 98262;
	#10 counter$count = 98263;
	#10 counter$count = 98264;
	#10 counter$count = 98265;
	#10 counter$count = 98266;
	#10 counter$count = 98267;
	#10 counter$count = 98268;
	#10 counter$count = 98269;
	#10 counter$count = 98270;
	#10 counter$count = 98271;
	#10 counter$count = 98272;
	#10 counter$count = 98273;
	#10 counter$count = 98274;
	#10 counter$count = 98275;
	#10 counter$count = 98276;
	#10 counter$count = 98277;
	#10 counter$count = 98278;
	#10 counter$count = 98279;
	#10 counter$count = 98280;
	#10 counter$count = 98281;
	#10 counter$count = 98282;
	#10 counter$count = 98283;
	#10 counter$count = 98284;
	#10 counter$count = 98285;
	#10 counter$count = 98286;
	#10 counter$count = 98287;
	#10 counter$count = 98288;
	#10 counter$count = 98289;
	#10 counter$count = 98290;
	#10 counter$count = 98291;
	#10 counter$count = 98292;
	#10 counter$count = 98293;
	#10 counter$count = 98294;
	#10 counter$count = 98295;
	#10 counter$count = 98296;
	#10 counter$count = 98297;
	#10 counter$count = 98298;
	#10 counter$count = 98299;
	#10 counter$count = 98300;
	#10 counter$count = 98301;
	#10 counter$count = 98302;
	#10 counter$count = 98303;
	#10 counter$count = 98304;
	#10 counter$count = 98305;
	#10 counter$count = 98306;
	#10 counter$count = 98307;
	#10 counter$count = 98308;
	#10 counter$count = 98309;
	#10 counter$count = 98310;
	#10 counter$count = 98311;
	#10 counter$count = 98312;
	#10 counter$count = 98313;
	#10 counter$count = 98314;
	#10 counter$count = 98315;
	#10 counter$count = 98316;
	#10 counter$count = 98317;
	#10 counter$count = 98318;
	#10 counter$count = 98319;
	#10 counter$count = 98320;
	#10 counter$count = 98321;
	#10 counter$count = 98322;
	#10 counter$count = 98323;
	#10 counter$count = 98324;
	#10 counter$count = 98325;
	#10 counter$count = 98326;
	#10 counter$count = 98327;
	#10 counter$count = 98328;
	#10 counter$count = 98329;
	#10 counter$count = 98330;
	#10 counter$count = 98331;
	#10 counter$count = 98332;
	#10 counter$count = 98333;
	#10 counter$count = 98334;
	#10 counter$count = 98335;
	#10 counter$count = 98336;
	#10 counter$count = 98337;
	#10 counter$count = 98338;
	#10 counter$count = 98339;
	#10 counter$count = 98340;
	#10 counter$count = 98341;
	#10 counter$count = 98342;
	#10 counter$count = 98343;
	#10 counter$count = 98344;
	#10 counter$count = 98345;
	#10 counter$count = 98346;
	#10 counter$count = 98347;
	#10 counter$count = 98348;
	#10 counter$count = 98349;
	#10 counter$count = 98350;
	#10 counter$count = 98351;
	#10 counter$count = 98352;
	#10 counter$count = 98353;
	#10 counter$count = 98354;
	#10 counter$count = 98355;
	#10 counter$count = 98356;
	#10 counter$count = 98357;
	#10 counter$count = 98358;
	#10 counter$count = 98359;
	#10 counter$count = 98360;
	#10 counter$count = 98361;
	#10 counter$count = 98362;
	#10 counter$count = 98363;
	#10 counter$count = 98364;
	#10 counter$count = 98365;
	#10 counter$count = 98366;
	#10 counter$count = 98367;
	#10 counter$count = 98368;
	#10 counter$count = 98369;
	#10 counter$count = 98370;
	#10 counter$count = 98371;
	#10 counter$count = 98372;
	#10 counter$count = 98373;
	#10 counter$count = 98374;
	#10 counter$count = 98375;
	#10 counter$count = 98376;
	#10 counter$count = 98377;
	#10 counter$count = 98378;
	#10 counter$count = 98379;
	#10 counter$count = 98380;
	#10 counter$count = 98381;
	#10 counter$count = 98382;
	#10 counter$count = 98383;
	#10 counter$count = 98384;
	#10 counter$count = 98385;
	#10 counter$count = 98386;
	#10 counter$count = 98387;
	#10 counter$count = 98388;
	#10 counter$count = 98389;
	#10 counter$count = 98390;
	#10 counter$count = 98391;
	#10 counter$count = 98392;
	#10 counter$count = 98393;
	#10 counter$count = 98394;
	#10 counter$count = 98395;
	#10 counter$count = 98396;
	#10 counter$count = 98397;
	#10 counter$count = 98398;
	#10 counter$count = 98399;
	#10 counter$count = 98400;
	#10 counter$count = 98401;
	#10 counter$count = 98402;
	#10 counter$count = 98403;
	#10 counter$count = 98404;
	#10 counter$count = 98405;
	#10 counter$count = 98406;
	#10 counter$count = 98407;
	#10 counter$count = 98408;
	#10 counter$count = 98409;
	#10 counter$count = 98410;
	#10 counter$count = 98411;
	#10 counter$count = 98412;
	#10 counter$count = 98413;
	#10 counter$count = 98414;
	#10 counter$count = 98415;
	#10 counter$count = 98416;
	#10 counter$count = 98417;
	#10 counter$count = 98418;
	#10 counter$count = 98419;
	#10 counter$count = 98420;
	#10 counter$count = 98421;
	#10 counter$count = 98422;
	#10 counter$count = 98423;
	#10 counter$count = 98424;
	#10 counter$count = 98425;
	#10 counter$count = 98426;
	#10 counter$count = 98427;
	#10 counter$count = 98428;
	#10 counter$count = 98429;
	#10 counter$count = 98430;
	#10 counter$count = 98431;
	#10 counter$count = 98432;
	#10 counter$count = 98433;
	#10 counter$count = 98434;
	#10 counter$count = 98435;
	#10 counter$count = 98436;
	#10 counter$count = 98437;
	#10 counter$count = 98438;
	#10 counter$count = 98439;
	#10 counter$count = 98440;
	#10 counter$count = 98441;
	#10 counter$count = 98442;
	#10 counter$count = 98443;
	#10 counter$count = 98444;
	#10 counter$count = 98445;
	#10 counter$count = 98446;
	#10 counter$count = 98447;
	#10 counter$count = 98448;
	#10 counter$count = 98449;
	#10 counter$count = 98450;
	#10 counter$count = 98451;
	#10 counter$count = 98452;
	#10 counter$count = 98453;
	#10 counter$count = 98454;
	#10 counter$count = 98455;
	#10 counter$count = 98456;
	#10 counter$count = 98457;
	#10 counter$count = 98458;
	#10 counter$count = 98459;
	#10 counter$count = 98460;
	#10 counter$count = 98461;
	#10 counter$count = 98462;
	#10 counter$count = 98463;
	#10 counter$count = 98464;
	#10 counter$count = 98465;
	#10 counter$count = 98466;
	#10 counter$count = 98467;
	#10 counter$count = 98468;
	#10 counter$count = 98469;
	#10 counter$count = 98470;
	#10 counter$count = 98471;
	#10 counter$count = 98472;
	#10 counter$count = 98473;
	#10 counter$count = 98474;
	#10 counter$count = 98475;
	#10 counter$count = 98476;
	#10 counter$count = 98477;
	#10 counter$count = 98478;
	#10 counter$count = 98479;
	#10 counter$count = 98480;
	#10 counter$count = 98481;
	#10 counter$count = 98482;
	#10 counter$count = 98483;
	#10 counter$count = 98484;
	#10 counter$count = 98485;
	#10 counter$count = 98486;
	#10 counter$count = 98487;
	#10 counter$count = 98488;
	#10 counter$count = 98489;
	#10 counter$count = 98490;
	#10 counter$count = 98491;
	#10 counter$count = 98492;
	#10 counter$count = 98493;
	#10 counter$count = 98494;
	#10 counter$count = 98495;
	#10 counter$count = 98496;
	#10 counter$count = 98497;
	#10 counter$count = 98498;
	#10 counter$count = 98499;
	#10 counter$count = 98500;
	#10 counter$count = 98501;
	#10 counter$count = 98502;
	#10 counter$count = 98503;
	#10 counter$count = 98504;
	#10 counter$count = 98505;
	#10 counter$count = 98506;
	#10 counter$count = 98507;
	#10 counter$count = 98508;
	#10 counter$count = 98509;
	#10 counter$count = 98510;
	#10 counter$count = 98511;
	#10 counter$count = 98512;
	#10 counter$count = 98513;
	#10 counter$count = 98514;
	#10 counter$count = 98515;
	#10 counter$count = 98516;
	#10 counter$count = 98517;
	#10 counter$count = 98518;
	#10 counter$count = 98519;
	#10 counter$count = 98520;
	#10 counter$count = 98521;
	#10 counter$count = 98522;
	#10 counter$count = 98523;
	#10 counter$count = 98524;
	#10 counter$count = 98525;
	#10 counter$count = 98526;
	#10 counter$count = 98527;
	#10 counter$count = 98528;
	#10 counter$count = 98529;
	#10 counter$count = 98530;
	#10 counter$count = 98531;
	#10 counter$count = 98532;
	#10 counter$count = 98533;
	#10 counter$count = 98534;
	#10 counter$count = 98535;
	#10 counter$count = 98536;
	#10 counter$count = 98537;
	#10 counter$count = 98538;
	#10 counter$count = 98539;
	#10 counter$count = 98540;
	#10 counter$count = 98541;
	#10 counter$count = 98542;
	#10 counter$count = 98543;
	#10 counter$count = 98544;
	#10 counter$count = 98545;
	#10 counter$count = 98546;
	#10 counter$count = 98547;
	#10 counter$count = 98548;
	#10 counter$count = 98549;
	#10 counter$count = 98550;
	#10 counter$count = 98551;
	#10 counter$count = 98552;
	#10 counter$count = 98553;
	#10 counter$count = 98554;
	#10 counter$count = 98555;
	#10 counter$count = 98556;
	#10 counter$count = 98557;
	#10 counter$count = 98558;
	#10 counter$count = 98559;
	#10 counter$count = 98560;
	#10 counter$count = 98561;
	#10 counter$count = 98562;
	#10 counter$count = 98563;
	#10 counter$count = 98564;
	#10 counter$count = 98565;
	#10 counter$count = 98566;
	#10 counter$count = 98567;
	#10 counter$count = 98568;
	#10 counter$count = 98569;
	#10 counter$count = 98570;
	#10 counter$count = 98571;
	#10 counter$count = 98572;
	#10 counter$count = 98573;
	#10 counter$count = 98574;
	#10 counter$count = 98575;
	#10 counter$count = 98576;
	#10 counter$count = 98577;
	#10 counter$count = 98578;
	#10 counter$count = 98579;
	#10 counter$count = 98580;
	#10 counter$count = 98581;
	#10 counter$count = 98582;
	#10 counter$count = 98583;
	#10 counter$count = 98584;
	#10 counter$count = 98585;
	#10 counter$count = 98586;
	#10 counter$count = 98587;
	#10 counter$count = 98588;
	#10 counter$count = 98589;
	#10 counter$count = 98590;
	#10 counter$count = 98591;
	#10 counter$count = 98592;
	#10 counter$count = 98593;
	#10 counter$count = 98594;
	#10 counter$count = 98595;
	#10 counter$count = 98596;
	#10 counter$count = 98597;
	#10 counter$count = 98598;
	#10 counter$count = 98599;
	#10 counter$count = 98600;
	#10 counter$count = 98601;
	#10 counter$count = 98602;
	#10 counter$count = 98603;
	#10 counter$count = 98604;
	#10 counter$count = 98605;
	#10 counter$count = 98606;
	#10 counter$count = 98607;
	#10 counter$count = 98608;
	#10 counter$count = 98609;
	#10 counter$count = 98610;
	#10 counter$count = 98611;
	#10 counter$count = 98612;
	#10 counter$count = 98613;
	#10 counter$count = 98614;
	#10 counter$count = 98615;
	#10 counter$count = 98616;
	#10 counter$count = 98617;
	#10 counter$count = 98618;
	#10 counter$count = 98619;
	#10 counter$count = 98620;
	#10 counter$count = 98621;
	#10 counter$count = 98622;
	#10 counter$count = 98623;
	#10 counter$count = 98624;
	#10 counter$count = 98625;
	#10 counter$count = 98626;
	#10 counter$count = 98627;
	#10 counter$count = 98628;
	#10 counter$count = 98629;
	#10 counter$count = 98630;
	#10 counter$count = 98631;
	#10 counter$count = 98632;
	#10 counter$count = 98633;
	#10 counter$count = 98634;
	#10 counter$count = 98635;
	#10 counter$count = 98636;
	#10 counter$count = 98637;
	#10 counter$count = 98638;
	#10 counter$count = 98639;
	#10 counter$count = 98640;
	#10 counter$count = 98641;
	#10 counter$count = 98642;
	#10 counter$count = 98643;
	#10 counter$count = 98644;
	#10 counter$count = 98645;
	#10 counter$count = 98646;
	#10 counter$count = 98647;
	#10 counter$count = 98648;
	#10 counter$count = 98649;
	#10 counter$count = 98650;
	#10 counter$count = 98651;
	#10 counter$count = 98652;
	#10 counter$count = 98653;
	#10 counter$count = 98654;
	#10 counter$count = 98655;
	#10 counter$count = 98656;
	#10 counter$count = 98657;
	#10 counter$count = 98658;
	#10 counter$count = 98659;
	#10 counter$count = 98660;
	#10 counter$count = 98661;
	#10 counter$count = 98662;
	#10 counter$count = 98663;
	#10 counter$count = 98664;
	#10 counter$count = 98665;
	#10 counter$count = 98666;
	#10 counter$count = 98667;
	#10 counter$count = 98668;
	#10 counter$count = 98669;
	#10 counter$count = 98670;
	#10 counter$count = 98671;
	#10 counter$count = 98672;
	#10 counter$count = 98673;
	#10 counter$count = 98674;
	#10 counter$count = 98675;
	#10 counter$count = 98676;
	#10 counter$count = 98677;
	#10 counter$count = 98678;
	#10 counter$count = 98679;
	#10 counter$count = 98680;
	#10 counter$count = 98681;
	#10 counter$count = 98682;
	#10 counter$count = 98683;
	#10 counter$count = 98684;
	#10 counter$count = 98685;
	#10 counter$count = 98686;
	#10 counter$count = 98687;
	#10 counter$count = 98688;
	#10 counter$count = 98689;
	#10 counter$count = 98690;
	#10 counter$count = 98691;
	#10 counter$count = 98692;
	#10 counter$count = 98693;
	#10 counter$count = 98694;
	#10 counter$count = 98695;
	#10 counter$count = 98696;
	#10 counter$count = 98697;
	#10 counter$count = 98698;
	#10 counter$count = 98699;
	#10 counter$count = 98700;
	#10 counter$count = 98701;
	#10 counter$count = 98702;
	#10 counter$count = 98703;
	#10 counter$count = 98704;
	#10 counter$count = 98705;
	#10 counter$count = 98706;
	#10 counter$count = 98707;
	#10 counter$count = 98708;
	#10 counter$count = 98709;
	#10 counter$count = 98710;
	#10 counter$count = 98711;
	#10 counter$count = 98712;
	#10 counter$count = 98713;
	#10 counter$count = 98714;
	#10 counter$count = 98715;
	#10 counter$count = 98716;
	#10 counter$count = 98717;
	#10 counter$count = 98718;
	#10 counter$count = 98719;
	#10 counter$count = 98720;
	#10 counter$count = 98721;
	#10 counter$count = 98722;
	#10 counter$count = 98723;
	#10 counter$count = 98724;
	#10 counter$count = 98725;
	#10 counter$count = 98726;
	#10 counter$count = 98727;
	#10 counter$count = 98728;
	#10 counter$count = 98729;
	#10 counter$count = 98730;
	#10 counter$count = 98731;
	#10 counter$count = 98732;
	#10 counter$count = 98733;
	#10 counter$count = 98734;
	#10 counter$count = 98735;
	#10 counter$count = 98736;
	#10 counter$count = 98737;
	#10 counter$count = 98738;
	#10 counter$count = 98739;
	#10 counter$count = 98740;
	#10 counter$count = 98741;
	#10 counter$count = 98742;
	#10 counter$count = 98743;
	#10 counter$count = 98744;
	#10 counter$count = 98745;
	#10 counter$count = 98746;
	#10 counter$count = 98747;
	#10 counter$count = 98748;
	#10 counter$count = 98749;
	#10 counter$count = 98750;
	#10 counter$count = 98751;
	#10 counter$count = 98752;
	#10 counter$count = 98753;
	#10 counter$count = 98754;
	#10 counter$count = 98755;
	#10 counter$count = 98756;
	#10 counter$count = 98757;
	#10 counter$count = 98758;
	#10 counter$count = 98759;
	#10 counter$count = 98760;
	#10 counter$count = 98761;
	#10 counter$count = 98762;
	#10 counter$count = 98763;
	#10 counter$count = 98764;
	#10 counter$count = 98765;
	#10 counter$count = 98766;
	#10 counter$count = 98767;
	#10 counter$count = 98768;
	#10 counter$count = 98769;
	#10 counter$count = 98770;
	#10 counter$count = 98771;
	#10 counter$count = 98772;
	#10 counter$count = 98773;
	#10 counter$count = 98774;
	#10 counter$count = 98775;
	#10 counter$count = 98776;
	#10 counter$count = 98777;
	#10 counter$count = 98778;
	#10 counter$count = 98779;
	#10 counter$count = 98780;
	#10 counter$count = 98781;
	#10 counter$count = 98782;
	#10 counter$count = 98783;
	#10 counter$count = 98784;
	#10 counter$count = 98785;
	#10 counter$count = 98786;
	#10 counter$count = 98787;
	#10 counter$count = 98788;
	#10 counter$count = 98789;
	#10 counter$count = 98790;
	#10 counter$count = 98791;
	#10 counter$count = 98792;
	#10 counter$count = 98793;
	#10 counter$count = 98794;
	#10 counter$count = 98795;
	#10 counter$count = 98796;
	#10 counter$count = 98797;
	#10 counter$count = 98798;
	#10 counter$count = 98799;
	#10 counter$count = 98800;
	#10 counter$count = 98801;
	#10 counter$count = 98802;
	#10 counter$count = 98803;
	#10 counter$count = 98804;
	#10 counter$count = 98805;
	#10 counter$count = 98806;
	#10 counter$count = 98807;
	#10 counter$count = 98808;
	#10 counter$count = 98809;
	#10 counter$count = 98810;
	#10 counter$count = 98811;
	#10 counter$count = 98812;
	#10 counter$count = 98813;
	#10 counter$count = 98814;
	#10 counter$count = 98815;
	#10 counter$count = 98816;
	#10 counter$count = 98817;
	#10 counter$count = 98818;
	#10 counter$count = 98819;
	#10 counter$count = 98820;
	#10 counter$count = 98821;
	#10 counter$count = 98822;
	#10 counter$count = 98823;
	#10 counter$count = 98824;
	#10 counter$count = 98825;
	#10 counter$count = 98826;
	#10 counter$count = 98827;
	#10 counter$count = 98828;
	#10 counter$count = 98829;
	#10 counter$count = 98830;
	#10 counter$count = 98831;
	#10 counter$count = 98832;
	#10 counter$count = 98833;
	#10 counter$count = 98834;
	#10 counter$count = 98835;
	#10 counter$count = 98836;
	#10 counter$count = 98837;
	#10 counter$count = 98838;
	#10 counter$count = 98839;
	#10 counter$count = 98840;
	#10 counter$count = 98841;
	#10 counter$count = 98842;
	#10 counter$count = 98843;
	#10 counter$count = 98844;
	#10 counter$count = 98845;
	#10 counter$count = 98846;
	#10 counter$count = 98847;
	#10 counter$count = 98848;
	#10 counter$count = 98849;
	#10 counter$count = 98850;
	#10 counter$count = 98851;
	#10 counter$count = 98852;
	#10 counter$count = 98853;
	#10 counter$count = 98854;
	#10 counter$count = 98855;
	#10 counter$count = 98856;
	#10 counter$count = 98857;
	#10 counter$count = 98858;
	#10 counter$count = 98859;
	#10 counter$count = 98860;
	#10 counter$count = 98861;
	#10 counter$count = 98862;
	#10 counter$count = 98863;
	#10 counter$count = 98864;
	#10 counter$count = 98865;
	#10 counter$count = 98866;
	#10 counter$count = 98867;
	#10 counter$count = 98868;
	#10 counter$count = 98869;
	#10 counter$count = 98870;
	#10 counter$count = 98871;
	#10 counter$count = 98872;
	#10 counter$count = 98873;
	#10 counter$count = 98874;
	#10 counter$count = 98875;
	#10 counter$count = 98876;
	#10 counter$count = 98877;
	#10 counter$count = 98878;
	#10 counter$count = 98879;
	#10 counter$count = 98880;
	#10 counter$count = 98881;
	#10 counter$count = 98882;
	#10 counter$count = 98883;
	#10 counter$count = 98884;
	#10 counter$count = 98885;
	#10 counter$count = 98886;
	#10 counter$count = 98887;
	#10 counter$count = 98888;
	#10 counter$count = 98889;
	#10 counter$count = 98890;
	#10 counter$count = 98891;
	#10 counter$count = 98892;
	#10 counter$count = 98893;
	#10 counter$count = 98894;
	#10 counter$count = 98895;
	#10 counter$count = 98896;
	#10 counter$count = 98897;
	#10 counter$count = 98898;
	#10 counter$count = 98899;
	#10 counter$count = 98900;
	#10 counter$count = 98901;
	#10 counter$count = 98902;
	#10 counter$count = 98903;
	#10 counter$count = 98904;
	#10 counter$count = 98905;
	#10 counter$count = 98906;
	#10 counter$count = 98907;
	#10 counter$count = 98908;
	#10 counter$count = 98909;
	#10 counter$count = 98910;
	#10 counter$count = 98911;
	#10 counter$count = 98912;
	#10 counter$count = 98913;
	#10 counter$count = 98914;
	#10 counter$count = 98915;
	#10 counter$count = 98916;
	#10 counter$count = 98917;
	#10 counter$count = 98918;
	#10 counter$count = 98919;
	#10 counter$count = 98920;
	#10 counter$count = 98921;
	#10 counter$count = 98922;
	#10 counter$count = 98923;
	#10 counter$count = 98924;
	#10 counter$count = 98925;
	#10 counter$count = 98926;
	#10 counter$count = 98927;
	#10 counter$count = 98928;
	#10 counter$count = 98929;
	#10 counter$count = 98930;
	#10 counter$count = 98931;
	#10 counter$count = 98932;
	#10 counter$count = 98933;
	#10 counter$count = 98934;
	#10 counter$count = 98935;
	#10 counter$count = 98936;
	#10 counter$count = 98937;
	#10 counter$count = 98938;
	#10 counter$count = 98939;
	#10 counter$count = 98940;
	#10 counter$count = 98941;
	#10 counter$count = 98942;
	#10 counter$count = 98943;
	#10 counter$count = 98944;
	#10 counter$count = 98945;
	#10 counter$count = 98946;
	#10 counter$count = 98947;
	#10 counter$count = 98948;
	#10 counter$count = 98949;
	#10 counter$count = 98950;
	#10 counter$count = 98951;
	#10 counter$count = 98952;
	#10 counter$count = 98953;
	#10 counter$count = 98954;
	#10 counter$count = 98955;
	#10 counter$count = 98956;
	#10 counter$count = 98957;
	#10 counter$count = 98958;
	#10 counter$count = 98959;
	#10 counter$count = 98960;
	#10 counter$count = 98961;
	#10 counter$count = 98962;
	#10 counter$count = 98963;
	#10 counter$count = 98964;
	#10 counter$count = 98965;
	#10 counter$count = 98966;
	#10 counter$count = 98967;
	#10 counter$count = 98968;
	#10 counter$count = 98969;
	#10 counter$count = 98970;
	#10 counter$count = 98971;
	#10 counter$count = 98972;
	#10 counter$count = 98973;
	#10 counter$count = 98974;
	#10 counter$count = 98975;
	#10 counter$count = 98976;
	#10 counter$count = 98977;
	#10 counter$count = 98978;
	#10 counter$count = 98979;
	#10 counter$count = 98980;
	#10 counter$count = 98981;
	#10 counter$count = 98982;
	#10 counter$count = 98983;
	#10 counter$count = 98984;
	#10 counter$count = 98985;
	#10 counter$count = 98986;
	#10 counter$count = 98987;
	#10 counter$count = 98988;
	#10 counter$count = 98989;
	#10 counter$count = 98990;
	#10 counter$count = 98991;
	#10 counter$count = 98992;
	#10 counter$count = 98993;
	#10 counter$count = 98994;
	#10 counter$count = 98995;
	#10 counter$count = 98996;
	#10 counter$count = 98997;
	#10 counter$count = 98998;
	#10 counter$count = 98999;
	#10 counter$count = 99000;
	#10 counter$count = 99001;
	#10 counter$count = 99002;
	#10 counter$count = 99003;
	#10 counter$count = 99004;
	#10 counter$count = 99005;
	#10 counter$count = 99006;
	#10 counter$count = 99007;
	#10 counter$count = 99008;
	#10 counter$count = 99009;
	#10 counter$count = 99010;
	#10 counter$count = 99011;
	#10 counter$count = 99012;
	#10 counter$count = 99013;
	#10 counter$count = 99014;
	#10 counter$count = 99015;
	#10 counter$count = 99016;
	#10 counter$count = 99017;
	#10 counter$count = 99018;
	#10 counter$count = 99019;
	#10 counter$count = 99020;
	#10 counter$count = 99021;
	#10 counter$count = 99022;
	#10 counter$count = 99023;
	#10 counter$count = 99024;
	#10 counter$count = 99025;
	#10 counter$count = 99026;
	#10 counter$count = 99027;
	#10 counter$count = 99028;
	#10 counter$count = 99029;
	#10 counter$count = 99030;
	#10 counter$count = 99031;
	#10 counter$count = 99032;
	#10 counter$count = 99033;
	#10 counter$count = 99034;
	#10 counter$count = 99035;
	#10 counter$count = 99036;
	#10 counter$count = 99037;
	#10 counter$count = 99038;
	#10 counter$count = 99039;
	#10 counter$count = 99040;
	#10 counter$count = 99041;
	#10 counter$count = 99042;
	#10 counter$count = 99043;
	#10 counter$count = 99044;
	#10 counter$count = 99045;
	#10 counter$count = 99046;
	#10 counter$count = 99047;
	#10 counter$count = 99048;
	#10 counter$count = 99049;
	#10 counter$count = 99050;
	#10 counter$count = 99051;
	#10 counter$count = 99052;
	#10 counter$count = 99053;
	#10 counter$count = 99054;
	#10 counter$count = 99055;
	#10 counter$count = 99056;
	#10 counter$count = 99057;
	#10 counter$count = 99058;
	#10 counter$count = 99059;
	#10 counter$count = 99060;
	#10 counter$count = 99061;
	#10 counter$count = 99062;
	#10 counter$count = 99063;
	#10 counter$count = 99064;
	#10 counter$count = 99065;
	#10 counter$count = 99066;
	#10 counter$count = 99067;
	#10 counter$count = 99068;
	#10 counter$count = 99069;
	#10 counter$count = 99070;
	#10 counter$count = 99071;
	#10 counter$count = 99072;
	#10 counter$count = 99073;
	#10 counter$count = 99074;
	#10 counter$count = 99075;
	#10 counter$count = 99076;
	#10 counter$count = 99077;
	#10 counter$count = 99078;
	#10 counter$count = 99079;
	#10 counter$count = 99080;
	#10 counter$count = 99081;
	#10 counter$count = 99082;
	#10 counter$count = 99083;
	#10 counter$count = 99084;
	#10 counter$count = 99085;
	#10 counter$count = 99086;
	#10 counter$count = 99087;
	#10 counter$count = 99088;
	#10 counter$count = 99089;
	#10 counter$count = 99090;
	#10 counter$count = 99091;
	#10 counter$count = 99092;
	#10 counter$count = 99093;
	#10 counter$count = 99094;
	#10 counter$count = 99095;
	#10 counter$count = 99096;
	#10 counter$count = 99097;
	#10 counter$count = 99098;
	#10 counter$count = 99099;
	#10 counter$count = 99100;
	#10 counter$count = 99101;
	#10 counter$count = 99102;
	#10 counter$count = 99103;
	#10 counter$count = 99104;
	#10 counter$count = 99105;
	#10 counter$count = 99106;
	#10 counter$count = 99107;
	#10 counter$count = 99108;
	#10 counter$count = 99109;
	#10 counter$count = 99110;
	#10 counter$count = 99111;
	#10 counter$count = 99112;
	#10 counter$count = 99113;
	#10 counter$count = 99114;
	#10 counter$count = 99115;
	#10 counter$count = 99116;
	#10 counter$count = 99117;
	#10 counter$count = 99118;
	#10 counter$count = 99119;
	#10 counter$count = 99120;
	#10 counter$count = 99121;
	#10 counter$count = 99122;
	#10 counter$count = 99123;
	#10 counter$count = 99124;
	#10 counter$count = 99125;
	#10 counter$count = 99126;
	#10 counter$count = 99127;
	#10 counter$count = 99128;
	#10 counter$count = 99129;
	#10 counter$count = 99130;
	#10 counter$count = 99131;
	#10 counter$count = 99132;
	#10 counter$count = 99133;
	#10 counter$count = 99134;
	#10 counter$count = 99135;
	#10 counter$count = 99136;
	#10 counter$count = 99137;
	#10 counter$count = 99138;
	#10 counter$count = 99139;
	#10 counter$count = 99140;
	#10 counter$count = 99141;
	#10 counter$count = 99142;
	#10 counter$count = 99143;
	#10 counter$count = 99144;
	#10 counter$count = 99145;
	#10 counter$count = 99146;
	#10 counter$count = 99147;
	#10 counter$count = 99148;
	#10 counter$count = 99149;
	#10 counter$count = 99150;
	#10 counter$count = 99151;
	#10 counter$count = 99152;
	#10 counter$count = 99153;
	#10 counter$count = 99154;
	#10 counter$count = 99155;
	#10 counter$count = 99156;
	#10 counter$count = 99157;
	#10 counter$count = 99158;
	#10 counter$count = 99159;
	#10 counter$count = 99160;
	#10 counter$count = 99161;
	#10 counter$count = 99162;
	#10 counter$count = 99163;
	#10 counter$count = 99164;
	#10 counter$count = 99165;
	#10 counter$count = 99166;
	#10 counter$count = 99167;
	#10 counter$count = 99168;
	#10 counter$count = 99169;
	#10 counter$count = 99170;
	#10 counter$count = 99171;
	#10 counter$count = 99172;
	#10 counter$count = 99173;
	#10 counter$count = 99174;
	#10 counter$count = 99175;
	#10 counter$count = 99176;
	#10 counter$count = 99177;
	#10 counter$count = 99178;
	#10 counter$count = 99179;
	#10 counter$count = 99180;
	#10 counter$count = 99181;
	#10 counter$count = 99182;
	#10 counter$count = 99183;
	#10 counter$count = 99184;
	#10 counter$count = 99185;
	#10 counter$count = 99186;
	#10 counter$count = 99187;
	#10 counter$count = 99188;
	#10 counter$count = 99189;
	#10 counter$count = 99190;
	#10 counter$count = 99191;
	#10 counter$count = 99192;
	#10 counter$count = 99193;
	#10 counter$count = 99194;
	#10 counter$count = 99195;
	#10 counter$count = 99196;
	#10 counter$count = 99197;
	#10 counter$count = 99198;
	#10 counter$count = 99199;
	#10 counter$count = 99200;
	#10 counter$count = 99201;
	#10 counter$count = 99202;
	#10 counter$count = 99203;
	#10 counter$count = 99204;
	#10 counter$count = 99205;
	#10 counter$count = 99206;
	#10 counter$count = 99207;
	#10 counter$count = 99208;
	#10 counter$count = 99209;
	#10 counter$count = 99210;
	#10 counter$count = 99211;
	#10 counter$count = 99212;
	#10 counter$count = 99213;
	#10 counter$count = 99214;
	#10 counter$count = 99215;
	#10 counter$count = 99216;
	#10 counter$count = 99217;
	#10 counter$count = 99218;
	#10 counter$count = 99219;
	#10 counter$count = 99220;
	#10 counter$count = 99221;
	#10 counter$count = 99222;
	#10 counter$count = 99223;
	#10 counter$count = 99224;
	#10 counter$count = 99225;
	#10 counter$count = 99226;
	#10 counter$count = 99227;
	#10 counter$count = 99228;
	#10 counter$count = 99229;
	#10 counter$count = 99230;
	#10 counter$count = 99231;
	#10 counter$count = 99232;
	#10 counter$count = 99233;
	#10 counter$count = 99234;
	#10 counter$count = 99235;
	#10 counter$count = 99236;
	#10 counter$count = 99237;
	#10 counter$count = 99238;
	#10 counter$count = 99239;
	#10 counter$count = 99240;
	#10 counter$count = 99241;
	#10 counter$count = 99242;
	#10 counter$count = 99243;
	#10 counter$count = 99244;
	#10 counter$count = 99245;
	#10 counter$count = 99246;
	#10 counter$count = 99247;
	#10 counter$count = 99248;
	#10 counter$count = 99249;
	#10 counter$count = 99250;
	#10 counter$count = 99251;
	#10 counter$count = 99252;
	#10 counter$count = 99253;
	#10 counter$count = 99254;
	#10 counter$count = 99255;
	#10 counter$count = 99256;
	#10 counter$count = 99257;
	#10 counter$count = 99258;
	#10 counter$count = 99259;
	#10 counter$count = 99260;
	#10 counter$count = 99261;
	#10 counter$count = 99262;
	#10 counter$count = 99263;
	#10 counter$count = 99264;
	#10 counter$count = 99265;
	#10 counter$count = 99266;
	#10 counter$count = 99267;
	#10 counter$count = 99268;
	#10 counter$count = 99269;
	#10 counter$count = 99270;
	#10 counter$count = 99271;
	#10 counter$count = 99272;
	#10 counter$count = 99273;
	#10 counter$count = 99274;
	#10 counter$count = 99275;
	#10 counter$count = 99276;
	#10 counter$count = 99277;
	#10 counter$count = 99278;
	#10 counter$count = 99279;
	#10 counter$count = 99280;
	#10 counter$count = 99281;
	#10 counter$count = 99282;
	#10 counter$count = 99283;
	#10 counter$count = 99284;
	#10 counter$count = 99285;
	#10 counter$count = 99286;
	#10 counter$count = 99287;
	#10 counter$count = 99288;
	#10 counter$count = 99289;
	#10 counter$count = 99290;
	#10 counter$count = 99291;
	#10 counter$count = 99292;
	#10 counter$count = 99293;
	#10 counter$count = 99294;
	#10 counter$count = 99295;
	#10 counter$count = 99296;
	#10 counter$count = 99297;
	#10 counter$count = 99298;
	#10 counter$count = 99299;
	#10 counter$count = 99300;
	#10 counter$count = 99301;
	#10 counter$count = 99302;
	#10 counter$count = 99303;
	#10 counter$count = 99304;
	#10 counter$count = 99305;
	#10 counter$count = 99306;
	#10 counter$count = 99307;
	#10 counter$count = 99308;
	#10 counter$count = 99309;
	#10 counter$count = 99310;
	#10 counter$count = 99311;
	#10 counter$count = 99312;
	#10 counter$count = 99313;
	#10 counter$count = 99314;
	#10 counter$count = 99315;
	#10 counter$count = 99316;
	#10 counter$count = 99317;
	#10 counter$count = 99318;
	#10 counter$count = 99319;
	#10 counter$count = 99320;
	#10 counter$count = 99321;
	#10 counter$count = 99322;
	#10 counter$count = 99323;
	#10 counter$count = 99324;
	#10 counter$count = 99325;
	#10 counter$count = 99326;
	#10 counter$count = 99327;
	#10 counter$count = 99328;
	#10 counter$count = 99329;
	#10 counter$count = 99330;
	#10 counter$count = 99331;
	#10 counter$count = 99332;
	#10 counter$count = 99333;
	#10 counter$count = 99334;
	#10 counter$count = 99335;
	#10 counter$count = 99336;
	#10 counter$count = 99337;
	#10 counter$count = 99338;
	#10 counter$count = 99339;
	#10 counter$count = 99340;
	#10 counter$count = 99341;
	#10 counter$count = 99342;
	#10 counter$count = 99343;
	#10 counter$count = 99344;
	#10 counter$count = 99345;
	#10 counter$count = 99346;
	#10 counter$count = 99347;
	#10 counter$count = 99348;
	#10 counter$count = 99349;
	#10 counter$count = 99350;
	#10 counter$count = 99351;
	#10 counter$count = 99352;
	#10 counter$count = 99353;
	#10 counter$count = 99354;
	#10 counter$count = 99355;
	#10 counter$count = 99356;
	#10 counter$count = 99357;
	#10 counter$count = 99358;
	#10 counter$count = 99359;
	#10 counter$count = 99360;
	#10 counter$count = 99361;
	#10 counter$count = 99362;
	#10 counter$count = 99363;
	#10 counter$count = 99364;
	#10 counter$count = 99365;
	#10 counter$count = 99366;
	#10 counter$count = 99367;
	#10 counter$count = 99368;
	#10 counter$count = 99369;
	#10 counter$count = 99370;
	#10 counter$count = 99371;
	#10 counter$count = 99372;
	#10 counter$count = 99373;
	#10 counter$count = 99374;
	#10 counter$count = 99375;
	#10 counter$count = 99376;
	#10 counter$count = 99377;
	#10 counter$count = 99378;
	#10 counter$count = 99379;
	#10 counter$count = 99380;
	#10 counter$count = 99381;
	#10 counter$count = 99382;
	#10 counter$count = 99383;
	#10 counter$count = 99384;
	#10 counter$count = 99385;
	#10 counter$count = 99386;
	#10 counter$count = 99387;
	#10 counter$count = 99388;
	#10 counter$count = 99389;
	#10 counter$count = 99390;
	#10 counter$count = 99391;
	#10 counter$count = 99392;
	#10 counter$count = 99393;
	#10 counter$count = 99394;
	#10 counter$count = 99395;
	#10 counter$count = 99396;
	#10 counter$count = 99397;
	#10 counter$count = 99398;
	#10 counter$count = 99399;
	#10 counter$count = 99400;
	#10 counter$count = 99401;
	#10 counter$count = 99402;
	#10 counter$count = 99403;
	#10 counter$count = 99404;
	#10 counter$count = 99405;
	#10 counter$count = 99406;
	#10 counter$count = 99407;
	#10 counter$count = 99408;
	#10 counter$count = 99409;
	#10 counter$count = 99410;
	#10 counter$count = 99411;
	#10 counter$count = 99412;
	#10 counter$count = 99413;
	#10 counter$count = 99414;
	#10 counter$count = 99415;
	#10 counter$count = 99416;
	#10 counter$count = 99417;
	#10 counter$count = 99418;
	#10 counter$count = 99419;
	#10 counter$count = 99420;
	#10 counter$count = 99421;
	#10 counter$count = 99422;
	#10 counter$count = 99423;
	#10 counter$count = 99424;
	#10 counter$count = 99425;
	#10 counter$count = 99426;
	#10 counter$count = 99427;
	#10 counter$count = 99428;
	#10 counter$count = 99429;
	#10 counter$count = 99430;
	#10 counter$count = 99431;
	#10 counter$count = 99432;
	#10 counter$count = 99433;
	#10 counter$count = 99434;
	#10 counter$count = 99435;
	#10 counter$count = 99436;
	#10 counter$count = 99437;
	#10 counter$count = 99438;
	#10 counter$count = 99439;
	#10 counter$count = 99440;
	#10 counter$count = 99441;
	#10 counter$count = 99442;
	#10 counter$count = 99443;
	#10 counter$count = 99444;
	#10 counter$count = 99445;
	#10 counter$count = 99446;
	#10 counter$count = 99447;
	#10 counter$count = 99448;
	#10 counter$count = 99449;
	#10 counter$count = 99450;
	#10 counter$count = 99451;
	#10 counter$count = 99452;
	#10 counter$count = 99453;
	#10 counter$count = 99454;
	#10 counter$count = 99455;
	#10 counter$count = 99456;
	#10 counter$count = 99457;
	#10 counter$count = 99458;
	#10 counter$count = 99459;
	#10 counter$count = 99460;
	#10 counter$count = 99461;
	#10 counter$count = 99462;
	#10 counter$count = 99463;
	#10 counter$count = 99464;
	#10 counter$count = 99465;
	#10 counter$count = 99466;
	#10 counter$count = 99467;
	#10 counter$count = 99468;
	#10 counter$count = 99469;
	#10 counter$count = 99470;
	#10 counter$count = 99471;
	#10 counter$count = 99472;
	#10 counter$count = 99473;
	#10 counter$count = 99474;
	#10 counter$count = 99475;
	#10 counter$count = 99476;
	#10 counter$count = 99477;
	#10 counter$count = 99478;
	#10 counter$count = 99479;
	#10 counter$count = 99480;
	#10 counter$count = 99481;
	#10 counter$count = 99482;
	#10 counter$count = 99483;
	#10 counter$count = 99484;
	#10 counter$count = 99485;
	#10 counter$count = 99486;
	#10 counter$count = 99487;
	#10 counter$count = 99488;
	#10 counter$count = 99489;
	#10 counter$count = 99490;
	#10 counter$count = 99491;
	#10 counter$count = 99492;
	#10 counter$count = 99493;
	#10 counter$count = 99494;
	#10 counter$count = 99495;
	#10 counter$count = 99496;
	#10 counter$count = 99497;
	#10 counter$count = 99498;
	#10 counter$count = 99499;
	#10 counter$count = 99500;
	#10 counter$count = 99501;
	#10 counter$count = 99502;
	#10 counter$count = 99503;
	#10 counter$count = 99504;
	#10 counter$count = 99505;
	#10 counter$count = 99506;
	#10 counter$count = 99507;
	#10 counter$count = 99508;
	#10 counter$count = 99509;
	#10 counter$count = 99510;
	#10 counter$count = 99511;
	#10 counter$count = 99512;
	#10 counter$count = 99513;
	#10 counter$count = 99514;
	#10 counter$count = 99515;
	#10 counter$count = 99516;
	#10 counter$count = 99517;
	#10 counter$count = 99518;
	#10 counter$count = 99519;
	#10 counter$count = 99520;
	#10 counter$count = 99521;
	#10 counter$count = 99522;
	#10 counter$count = 99523;
	#10 counter$count = 99524;
	#10 counter$count = 99525;
	#10 counter$count = 99526;
	#10 counter$count = 99527;
	#10 counter$count = 99528;
	#10 counter$count = 99529;
	#10 counter$count = 99530;
	#10 counter$count = 99531;
	#10 counter$count = 99532;
	#10 counter$count = 99533;
	#10 counter$count = 99534;
	#10 counter$count = 99535;
	#10 counter$count = 99536;
	#10 counter$count = 99537;
	#10 counter$count = 99538;
	#10 counter$count = 99539;
	#10 counter$count = 99540;
	#10 counter$count = 99541;
	#10 counter$count = 99542;
	#10 counter$count = 99543;
	#10 counter$count = 99544;
	#10 counter$count = 99545;
	#10 counter$count = 99546;
	#10 counter$count = 99547;
	#10 counter$count = 99548;
	#10 counter$count = 99549;
	#10 counter$count = 99550;
	#10 counter$count = 99551;
	#10 counter$count = 99552;
	#10 counter$count = 99553;
	#10 counter$count = 99554;
	#10 counter$count = 99555;
	#10 counter$count = 99556;
	#10 counter$count = 99557;
	#10 counter$count = 99558;
	#10 counter$count = 99559;
	#10 counter$count = 99560;
	#10 counter$count = 99561;
	#10 counter$count = 99562;
	#10 counter$count = 99563;
	#10 counter$count = 99564;
	#10 counter$count = 99565;
	#10 counter$count = 99566;
	#10 counter$count = 99567;
	#10 counter$count = 99568;
	#10 counter$count = 99569;
	#10 counter$count = 99570;
	#10 counter$count = 99571;
	#10 counter$count = 99572;
	#10 counter$count = 99573;
	#10 counter$count = 99574;
	#10 counter$count = 99575;
	#10 counter$count = 99576;
	#10 counter$count = 99577;
	#10 counter$count = 99578;
	#10 counter$count = 99579;
	#10 counter$count = 99580;
	#10 counter$count = 99581;
	#10 counter$count = 99582;
	#10 counter$count = 99583;
	#10 counter$count = 99584;
	#10 counter$count = 99585;
	#10 counter$count = 99586;
	#10 counter$count = 99587;
	#10 counter$count = 99588;
	#10 counter$count = 99589;
	#10 counter$count = 99590;
	#10 counter$count = 99591;
	#10 counter$count = 99592;
	#10 counter$count = 99593;
	#10 counter$count = 99594;
	#10 counter$count = 99595;
	#10 counter$count = 99596;
	#10 counter$count = 99597;
	#10 counter$count = 99598;
	#10 counter$count = 99599;
	#10 counter$count = 99600;
	#10 counter$count = 99601;
	#10 counter$count = 99602;
	#10 counter$count = 99603;
	#10 counter$count = 99604;
	#10 counter$count = 99605;
	#10 counter$count = 99606;
	#10 counter$count = 99607;
	#10 counter$count = 99608;
	#10 counter$count = 99609;
	#10 counter$count = 99610;
	#10 counter$count = 99611;
	#10 counter$count = 99612;
	#10 counter$count = 99613;
	#10 counter$count = 99614;
	#10 counter$count = 99615;
	#10 counter$count = 99616;
	#10 counter$count = 99617;
	#10 counter$count = 99618;
	#10 counter$count = 99619;
	#10 counter$count = 99620;
	#10 counter$count = 99621;
	#10 counter$count = 99622;
	#10 counter$count = 99623;
	#10 counter$count = 99624;
	#10 counter$count = 99625;
	#10 counter$count = 99626;
	#10 counter$count = 99627;
	#10 counter$count = 99628;
	#10 counter$count = 99629;
	#10 counter$count = 99630;
	#10 counter$count = 99631;
	#10 counter$count = 99632;
	#10 counter$count = 99633;
	#10 counter$count = 99634;
	#10 counter$count = 99635;
	#10 counter$count = 99636;
	#10 counter$count = 99637;
	#10 counter$count = 99638;
	#10 counter$count = 99639;
	#10 counter$count = 99640;
	#10 counter$count = 99641;
	#10 counter$count = 99642;
	#10 counter$count = 99643;
	#10 counter$count = 99644;
	#10 counter$count = 99645;
	#10 counter$count = 99646;
	#10 counter$count = 99647;
	#10 counter$count = 99648;
	#10 counter$count = 99649;
	#10 counter$count = 99650;
	#10 counter$count = 99651;
	#10 counter$count = 99652;
	#10 counter$count = 99653;
	#10 counter$count = 99654;
	#10 counter$count = 99655;
	#10 counter$count = 99656;
	#10 counter$count = 99657;
	#10 counter$count = 99658;
	#10 counter$count = 99659;
	#10 counter$count = 99660;
	#10 counter$count = 99661;
	#10 counter$count = 99662;
	#10 counter$count = 99663;
	#10 counter$count = 99664;
	#10 counter$count = 99665;
	#10 counter$count = 99666;
	#10 counter$count = 99667;
	#10 counter$count = 99668;
	#10 counter$count = 99669;
	#10 counter$count = 99670;
	#10 counter$count = 99671;
	#10 counter$count = 99672;
	#10 counter$count = 99673;
	#10 counter$count = 99674;
	#10 counter$count = 99675;
	#10 counter$count = 99676;
	#10 counter$count = 99677;
	#10 counter$count = 99678;
	#10 counter$count = 99679;
	#10 counter$count = 99680;
	#10 counter$count = 99681;
	#10 counter$count = 99682;
	#10 counter$count = 99683;
	#10 counter$count = 99684;
	#10 counter$count = 99685;
	#10 counter$count = 99686;
	#10 counter$count = 99687;
	#10 counter$count = 99688;
	#10 counter$count = 99689;
	#10 counter$count = 99690;
	#10 counter$count = 99691;
	#10 counter$count = 99692;
	#10 counter$count = 99693;
	#10 counter$count = 99694;
	#10 counter$count = 99695;
	#10 counter$count = 99696;
	#10 counter$count = 99697;
	#10 counter$count = 99698;
	#10 counter$count = 99699;
	#10 counter$count = 99700;
	#10 counter$count = 99701;
	#10 counter$count = 99702;
	#10 counter$count = 99703;
	#10 counter$count = 99704;
	#10 counter$count = 99705;
	#10 counter$count = 99706;
	#10 counter$count = 99707;
	#10 counter$count = 99708;
	#10 counter$count = 99709;
	#10 counter$count = 99710;
	#10 counter$count = 99711;
	#10 counter$count = 99712;
	#10 counter$count = 99713;
	#10 counter$count = 99714;
	#10 counter$count = 99715;
	#10 counter$count = 99716;
	#10 counter$count = 99717;
	#10 counter$count = 99718;
	#10 counter$count = 99719;
	#10 counter$count = 99720;
	#10 counter$count = 99721;
	#10 counter$count = 99722;
	#10 counter$count = 99723;
	#10 counter$count = 99724;
	#10 counter$count = 99725;
	#10 counter$count = 99726;
	#10 counter$count = 99727;
	#10 counter$count = 99728;
	#10 counter$count = 99729;
	#10 counter$count = 99730;
	#10 counter$count = 99731;
	#10 counter$count = 99732;
	#10 counter$count = 99733;
	#10 counter$count = 99734;
	#10 counter$count = 99735;
	#10 counter$count = 99736;
	#10 counter$count = 99737;
	#10 counter$count = 99738;
	#10 counter$count = 99739;
	#10 counter$count = 99740;
	#10 counter$count = 99741;
	#10 counter$count = 99742;
	#10 counter$count = 99743;
	#10 counter$count = 99744;
	#10 counter$count = 99745;
	#10 counter$count = 99746;
	#10 counter$count = 99747;
	#10 counter$count = 99748;
	#10 counter$count = 99749;
	#10 counter$count = 99750;
	#10 counter$count = 99751;
	#10 counter$count = 99752;
	#10 counter$count = 99753;
	#10 counter$count = 99754;
	#10 counter$count = 99755;
	#10 counter$count = 99756;
	#10 counter$count = 99757;
	#10 counter$count = 99758;
	#10 counter$count = 99759;
	#10 counter$count = 99760;
	#10 counter$count = 99761;
	#10 counter$count = 99762;
	#10 counter$count = 99763;
	#10 counter$count = 99764;
	#10 counter$count = 99765;
	#10 counter$count = 99766;
	#10 counter$count = 99767;
	#10 counter$count = 99768;
	#10 counter$count = 99769;
	#10 counter$count = 99770;
	#10 counter$count = 99771;
	#10 counter$count = 99772;
	#10 counter$count = 99773;
	#10 counter$count = 99774;
	#10 counter$count = 99775;
	#10 counter$count = 99776;
	#10 counter$count = 99777;
	#10 counter$count = 99778;
	#10 counter$count = 99779;
	#10 counter$count = 99780;
	#10 counter$count = 99781;
	#10 counter$count = 99782;
	#10 counter$count = 99783;
	#10 counter$count = 99784;
	#10 counter$count = 99785;
	#10 counter$count = 99786;
	#10 counter$count = 99787;
	#10 counter$count = 99788;
	#10 counter$count = 99789;
	#10 counter$count = 99790;
	#10 counter$count = 99791;
	#10 counter$count = 99792;
	#10 counter$count = 99793;
	#10 counter$count = 99794;
	#10 counter$count = 99795;
	#10 counter$count = 99796;
	#10 counter$count = 99797;
	#10 counter$count = 99798;
	#10 counter$count = 99799;
	#10 counter$count = 99800;
	#10 counter$count = 99801;
	#10 counter$count = 99802;
	#10 counter$count = 99803;
	#10 counter$count = 99804;
	#10 counter$count = 99805;
	#10 counter$count = 99806;
	#10 counter$count = 99807;
	#10 counter$count = 99808;
	#10 counter$count = 99809;
	#10 counter$count = 99810;
	#10 counter$count = 99811;
	#10 counter$count = 99812;
	#10 counter$count = 99813;
	#10 counter$count = 99814;
	#10 counter$count = 99815;
	#10 counter$count = 99816;
	#10 counter$count = 99817;
	#10 counter$count = 99818;
	#10 counter$count = 99819;
	#10 counter$count = 99820;
	#10 counter$count = 99821;
	#10 counter$count = 99822;
	#10 counter$count = 99823;
	#10 counter$count = 99824;
	#10 counter$count = 99825;
	#10 counter$count = 99826;
	#10 counter$count = 99827;
	#10 counter$count = 99828;
	#10 counter$count = 99829;
	#10 counter$count = 99830;
	#10 counter$count = 99831;
	#10 counter$count = 99832;
	#10 counter$count = 99833;
	#10 counter$count = 99834;
	#10 counter$count = 99835;
	#10 counter$count = 99836;
	#10 counter$count = 99837;
	#10 counter$count = 99838;
	#10 counter$count = 99839;
	#10 counter$count = 99840;
	#10 counter$count = 99841;
	#10 counter$count = 99842;
	#10 counter$count = 99843;
	#10 counter$count = 99844;
	#10 counter$count = 99845;
	#10 counter$count = 99846;
	#10 counter$count = 99847;
	#10 counter$count = 99848;
	#10 counter$count = 99849;
	#10 counter$count = 99850;
	#10 counter$count = 99851;
	#10 counter$count = 99852;
	#10 counter$count = 99853;
	#10 counter$count = 99854;
	#10 counter$count = 99855;
	#10 counter$count = 99856;
	#10 counter$count = 99857;
	#10 counter$count = 99858;
	#10 counter$count = 99859;
	#10 counter$count = 99860;
	#10 counter$count = 99861;
	#10 counter$count = 99862;
	#10 counter$count = 99863;
	#10 counter$count = 99864;
	#10 counter$count = 99865;
	#10 counter$count = 99866;
	#10 counter$count = 99867;
	#10 counter$count = 99868;
	#10 counter$count = 99869;
	#10 counter$count = 99870;
	#10 counter$count = 99871;
	#10 counter$count = 99872;
	#10 counter$count = 99873;
	#10 counter$count = 99874;
	#10 counter$count = 99875;
	#10 counter$count = 99876;
	#10 counter$count = 99877;
	#10 counter$count = 99878;
	#10 counter$count = 99879;
	#10 counter$count = 99880;
	#10 counter$count = 99881;
	#10 counter$count = 99882;
	#10 counter$count = 99883;
	#10 counter$count = 99884;
	#10 counter$count = 99885;
	#10 counter$count = 99886;
	#10 counter$count = 99887;
	#10 counter$count = 99888;
	#10 counter$count = 99889;
	#10 counter$count = 99890;
	#10 counter$count = 99891;
	#10 counter$count = 99892;
	#10 counter$count = 99893;
	#10 counter$count = 99894;
	#10 counter$count = 99895;
	#10 counter$count = 99896;
	#10 counter$count = 99897;
	#10 counter$count = 99898;
	#10 counter$count = 99899;
	#10 counter$count = 99900;
	#10 counter$count = 99901;
	#10 counter$count = 99902;
	#10 counter$count = 99903;
	#10 counter$count = 99904;
	#10 counter$count = 99905;
	#10 counter$count = 99906;
	#10 counter$count = 99907;
	#10 counter$count = 99908;
	#10 counter$count = 99909;
	#10 counter$count = 99910;
	#10 counter$count = 99911;
	#10 counter$count = 99912;
	#10 counter$count = 99913;
	#10 counter$count = 99914;
	#10 counter$count = 99915;
	#10 counter$count = 99916;
	#10 counter$count = 99917;
	#10 counter$count = 99918;
	#10 counter$count = 99919;
	#10 counter$count = 99920;
	#10 counter$count = 99921;
	#10 counter$count = 99922;
	#10 counter$count = 99923;
	#10 counter$count = 99924;
	#10 counter$count = 99925;
	#10 counter$count = 99926;
	#10 counter$count = 99927;
	#10 counter$count = 99928;
	#10 counter$count = 99929;
	#10 counter$count = 99930;
	#10 counter$count = 99931;
	#10 counter$count = 99932;
	#10 counter$count = 99933;
	#10 counter$count = 99934;
	#10 counter$count = 99935;
	#10 counter$count = 99936;
	#10 counter$count = 99937;
	#10 counter$count = 99938;
	#10 counter$count = 99939;
	#10 counter$count = 99940;
	#10 counter$count = 99941;
	#10 counter$count = 99942;
	#10 counter$count = 99943;
	#10 counter$count = 99944;
	#10 counter$count = 99945;
	#10 counter$count = 99946;
	#10 counter$count = 99947;
	#10 counter$count = 99948;
	#10 counter$count = 99949;
	#10 counter$count = 99950;
	#10 counter$count = 99951;
	#10 counter$count = 99952;
	#10 counter$count = 99953;
	#10 counter$count = 99954;
	#10 counter$count = 99955;
	#10 counter$count = 99956;
	#10 counter$count = 99957;
	#10 counter$count = 99958;
	#10 counter$count = 99959;
	#10 counter$count = 99960;
	#10 counter$count = 99961;
	#10 counter$count = 99962;
	#10 counter$count = 99963;
	#10 counter$count = 99964;
	#10 counter$count = 99965;
	#10 counter$count = 99966;
	#10 counter$count = 99967;
	#10 counter$count = 99968;
	#10 counter$count = 99969;
	#10 counter$count = 99970;
	#10 counter$count = 99971;
	#10 counter$count = 99972;
	#10 counter$count = 99973;
	#10 counter$count = 99974;
	#10 counter$count = 99975;
	#10 counter$count = 99976;
	#10 counter$count = 99977;
	#10 counter$count = 99978;
	#10 counter$count = 99979;
	#10 counter$count = 99980;
	#10 counter$count = 99981;
	#10 counter$count = 99982;
	#10 counter$count = 99983;
	#10 counter$count = 99984;
	#10 counter$count = 99985;
	#10 counter$count = 99986;
	#10 counter$count = 99987;
	#10 counter$count = 99988;
	#10 counter$count = 99989;
	#10 counter$count = 99990;
	#10 counter$count = 99991;
	#10 counter$count = 99992;
	#10 counter$count = 99993;
	#10 counter$count = 99994;
	#10 counter$count = 99995;
	#10 counter$count = 99996;
	#10 counter$count = 99997;
	#10 counter$count = 99998;
	#10 counter$count = 99999;
	#10 counter$count = 100000;
	#10 counter$count = 100001;
end
 // port: counter$overflow
initial begin
	#0 counter$overflow = 0;
end
 // for en_regs 

initial begin
	#1000020 $finish;
end
initial begin
	$dumpfile("tb$top.vcd");
	$dumpvars(0, testbench);
end
endmodule

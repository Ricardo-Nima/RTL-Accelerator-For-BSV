`timescale 1ns/1ns
module testbench();
 reg CLK, RST_N;
 reg [2 : 0] spi_writer$spi;
 reg [7 : 0] spi_writer$hook_write_data;
 mkDecCounter U1(.CLK(CLK), 
		.RST_N(RST_N), 
		.spi_writer$spi(spi_writer$spi), 
		.spi_writer$hook_write_data(spi_writer$hook_write_data), 
		.count(), 
		.RDY_count(), 
		.overflow(), 
		.RDY_overflow());
always begin
	#5 CLK = ~CLK;
end
initial begin
	RST_N = 0;
	#1 CLK = 1;
	#1 RST_N = 1;
end
 // port: spi_writer$spi
initial begin
	#0 spi_writer$spi = 0;
	#10 spi_writer$spi = 7;
	#20 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 7;
	#30 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#10 spi_writer$spi = 0;
	#10 spi_writer$spi = 2;
	#10 spi_writer$spi = 1;
	#10 spi_writer$spi = 3;
	#20 spi_writer$spi = 7;
end
 // port: spi_writer$hook_write_data
initial begin
	#0 spi_writer$hook_write_data = 170;
	#10 spi_writer$hook_write_data = 0;
	#220 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
	#210 spi_writer$hook_write_data = 162;
	#210 spi_writer$hook_write_data = 183;
	#210 spi_writer$hook_write_data = 204;
	#210 spi_writer$hook_write_data = 225;
	#210 spi_writer$hook_write_data = 246;
	#210 spi_writer$hook_write_data = 11;
	#210 spi_writer$hook_write_data = 32;
	#210 spi_writer$hook_write_data = 53;
	#210 spi_writer$hook_write_data = 74;
	#210 spi_writer$hook_write_data = 95;
	#210 spi_writer$hook_write_data = 116;
	#210 spi_writer$hook_write_data = 137;
	#210 spi_writer$hook_write_data = 158;
	#210 spi_writer$hook_write_data = 179;
	#210 spi_writer$hook_write_data = 200;
	#210 spi_writer$hook_write_data = 221;
	#210 spi_writer$hook_write_data = 242;
	#210 spi_writer$hook_write_data = 7;
	#210 spi_writer$hook_write_data = 28;
	#210 spi_writer$hook_write_data = 49;
	#210 spi_writer$hook_write_data = 70;
	#210 spi_writer$hook_write_data = 91;
	#210 spi_writer$hook_write_data = 112;
	#210 spi_writer$hook_write_data = 133;
	#210 spi_writer$hook_write_data = 154;
	#210 spi_writer$hook_write_data = 175;
	#210 spi_writer$hook_write_data = 196;
	#210 spi_writer$hook_write_data = 217;
	#210 spi_writer$hook_write_data = 238;
	#210 spi_writer$hook_write_data = 3;
	#210 spi_writer$hook_write_data = 24;
	#210 spi_writer$hook_write_data = 45;
	#210 spi_writer$hook_write_data = 66;
	#210 spi_writer$hook_write_data = 87;
	#210 spi_writer$hook_write_data = 108;
	#210 spi_writer$hook_write_data = 129;
	#210 spi_writer$hook_write_data = 150;
	#210 spi_writer$hook_write_data = 171;
	#210 spi_writer$hook_write_data = 192;
	#210 spi_writer$hook_write_data = 213;
	#210 spi_writer$hook_write_data = 234;
	#210 spi_writer$hook_write_data = 255;
	#210 spi_writer$hook_write_data = 20;
	#210 spi_writer$hook_write_data = 41;
	#210 spi_writer$hook_write_data = 62;
	#210 spi_writer$hook_write_data = 83;
	#210 spi_writer$hook_write_data = 104;
	#210 spi_writer$hook_write_data = 125;
	#210 spi_writer$hook_write_data = 146;
	#210 spi_writer$hook_write_data = 167;
	#210 spi_writer$hook_write_data = 188;
	#210 spi_writer$hook_write_data = 209;
	#210 spi_writer$hook_write_data = 230;
	#210 spi_writer$hook_write_data = 251;
	#210 spi_writer$hook_write_data = 16;
	#210 spi_writer$hook_write_data = 37;
	#210 spi_writer$hook_write_data = 58;
	#210 spi_writer$hook_write_data = 79;
	#210 spi_writer$hook_write_data = 100;
	#210 spi_writer$hook_write_data = 121;
	#210 spi_writer$hook_write_data = 142;
	#210 spi_writer$hook_write_data = 163;
	#210 spi_writer$hook_write_data = 184;
	#210 spi_writer$hook_write_data = 205;
	#210 spi_writer$hook_write_data = 226;
	#210 spi_writer$hook_write_data = 247;
	#210 spi_writer$hook_write_data = 12;
	#210 spi_writer$hook_write_data = 33;
	#210 spi_writer$hook_write_data = 54;
	#210 spi_writer$hook_write_data = 75;
	#210 spi_writer$hook_write_data = 96;
	#210 spi_writer$hook_write_data = 117;
	#210 spi_writer$hook_write_data = 138;
	#210 spi_writer$hook_write_data = 159;
	#210 spi_writer$hook_write_data = 180;
	#210 spi_writer$hook_write_data = 201;
	#210 spi_writer$hook_write_data = 222;
	#210 spi_writer$hook_write_data = 243;
	#210 spi_writer$hook_write_data = 8;
	#210 spi_writer$hook_write_data = 29;
	#210 spi_writer$hook_write_data = 50;
	#210 spi_writer$hook_write_data = 71;
	#210 spi_writer$hook_write_data = 92;
	#210 spi_writer$hook_write_data = 113;
	#210 spi_writer$hook_write_data = 134;
	#210 spi_writer$hook_write_data = 155;
	#210 spi_writer$hook_write_data = 176;
	#210 spi_writer$hook_write_data = 197;
	#210 spi_writer$hook_write_data = 218;
	#210 spi_writer$hook_write_data = 239;
	#210 spi_writer$hook_write_data = 4;
	#210 spi_writer$hook_write_data = 25;
	#210 spi_writer$hook_write_data = 46;
	#210 spi_writer$hook_write_data = 67;
	#210 spi_writer$hook_write_data = 88;
	#210 spi_writer$hook_write_data = 109;
	#210 spi_writer$hook_write_data = 130;
	#210 spi_writer$hook_write_data = 151;
	#210 spi_writer$hook_write_data = 172;
	#210 spi_writer$hook_write_data = 193;
	#210 spi_writer$hook_write_data = 214;
	#210 spi_writer$hook_write_data = 235;
	#210 spi_writer$hook_write_data = 0;
	#210 spi_writer$hook_write_data = 21;
	#210 spi_writer$hook_write_data = 42;
	#210 spi_writer$hook_write_data = 63;
	#210 spi_writer$hook_write_data = 84;
	#210 spi_writer$hook_write_data = 105;
	#210 spi_writer$hook_write_data = 126;
	#210 spi_writer$hook_write_data = 147;
	#210 spi_writer$hook_write_data = 168;
	#210 spi_writer$hook_write_data = 189;
	#210 spi_writer$hook_write_data = 210;
	#210 spi_writer$hook_write_data = 231;
	#210 spi_writer$hook_write_data = 252;
	#210 spi_writer$hook_write_data = 17;
	#210 spi_writer$hook_write_data = 38;
	#210 spi_writer$hook_write_data = 59;
	#210 spi_writer$hook_write_data = 80;
	#210 spi_writer$hook_write_data = 101;
	#210 spi_writer$hook_write_data = 122;
	#210 spi_writer$hook_write_data = 143;
	#210 spi_writer$hook_write_data = 164;
	#210 spi_writer$hook_write_data = 185;
	#210 spi_writer$hook_write_data = 206;
	#210 spi_writer$hook_write_data = 227;
	#210 spi_writer$hook_write_data = 248;
	#210 spi_writer$hook_write_data = 13;
	#210 spi_writer$hook_write_data = 34;
	#210 spi_writer$hook_write_data = 55;
	#210 spi_writer$hook_write_data = 76;
	#210 spi_writer$hook_write_data = 97;
	#210 spi_writer$hook_write_data = 118;
	#210 spi_writer$hook_write_data = 139;
	#210 spi_writer$hook_write_data = 160;
	#210 spi_writer$hook_write_data = 181;
	#210 spi_writer$hook_write_data = 202;
	#210 spi_writer$hook_write_data = 223;
	#210 spi_writer$hook_write_data = 244;
	#210 spi_writer$hook_write_data = 9;
	#210 spi_writer$hook_write_data = 30;
	#210 spi_writer$hook_write_data = 51;
	#210 spi_writer$hook_write_data = 72;
	#210 spi_writer$hook_write_data = 93;
	#210 spi_writer$hook_write_data = 114;
	#210 spi_writer$hook_write_data = 135;
	#210 spi_writer$hook_write_data = 156;
	#210 spi_writer$hook_write_data = 177;
	#210 spi_writer$hook_write_data = 198;
	#210 spi_writer$hook_write_data = 219;
	#210 spi_writer$hook_write_data = 240;
	#210 spi_writer$hook_write_data = 5;
	#210 spi_writer$hook_write_data = 26;
	#210 spi_writer$hook_write_data = 47;
	#210 spi_writer$hook_write_data = 68;
	#210 spi_writer$hook_write_data = 89;
	#210 spi_writer$hook_write_data = 110;
	#210 spi_writer$hook_write_data = 131;
	#210 spi_writer$hook_write_data = 152;
	#210 spi_writer$hook_write_data = 173;
	#210 spi_writer$hook_write_data = 194;
	#210 spi_writer$hook_write_data = 215;
	#210 spi_writer$hook_write_data = 236;
	#210 spi_writer$hook_write_data = 1;
	#210 spi_writer$hook_write_data = 22;
	#210 spi_writer$hook_write_data = 43;
	#210 spi_writer$hook_write_data = 64;
	#210 spi_writer$hook_write_data = 85;
	#210 spi_writer$hook_write_data = 106;
	#210 spi_writer$hook_write_data = 127;
	#210 spi_writer$hook_write_data = 148;
	#210 spi_writer$hook_write_data = 169;
	#210 spi_writer$hook_write_data = 190;
	#210 spi_writer$hook_write_data = 211;
	#210 spi_writer$hook_write_data = 232;
	#210 spi_writer$hook_write_data = 253;
	#210 spi_writer$hook_write_data = 18;
	#210 spi_writer$hook_write_data = 39;
	#210 spi_writer$hook_write_data = 60;
	#210 spi_writer$hook_write_data = 81;
	#210 spi_writer$hook_write_data = 102;
	#210 spi_writer$hook_write_data = 123;
	#210 spi_writer$hook_write_data = 144;
	#210 spi_writer$hook_write_data = 165;
	#210 spi_writer$hook_write_data = 186;
	#210 spi_writer$hook_write_data = 207;
	#210 spi_writer$hook_write_data = 228;
	#210 spi_writer$hook_write_data = 249;
	#210 spi_writer$hook_write_data = 14;
	#210 spi_writer$hook_write_data = 35;
	#210 spi_writer$hook_write_data = 56;
	#210 spi_writer$hook_write_data = 77;
	#210 spi_writer$hook_write_data = 98;
	#210 spi_writer$hook_write_data = 119;
	#210 spi_writer$hook_write_data = 140;
	#210 spi_writer$hook_write_data = 161;
	#210 spi_writer$hook_write_data = 182;
	#210 spi_writer$hook_write_data = 203;
	#210 spi_writer$hook_write_data = 224;
	#210 spi_writer$hook_write_data = 245;
	#210 spi_writer$hook_write_data = 10;
	#210 spi_writer$hook_write_data = 31;
	#210 spi_writer$hook_write_data = 52;
	#210 spi_writer$hook_write_data = 73;
	#210 spi_writer$hook_write_data = 94;
	#210 spi_writer$hook_write_data = 115;
	#210 spi_writer$hook_write_data = 136;
	#210 spi_writer$hook_write_data = 157;
	#210 spi_writer$hook_write_data = 178;
	#210 spi_writer$hook_write_data = 199;
	#210 spi_writer$hook_write_data = 220;
	#210 spi_writer$hook_write_data = 241;
	#210 spi_writer$hook_write_data = 6;
	#210 spi_writer$hook_write_data = 27;
	#210 spi_writer$hook_write_data = 48;
	#210 spi_writer$hook_write_data = 69;
	#210 spi_writer$hook_write_data = 90;
	#210 spi_writer$hook_write_data = 111;
	#210 spi_writer$hook_write_data = 132;
	#210 spi_writer$hook_write_data = 153;
	#210 spi_writer$hook_write_data = 174;
	#210 spi_writer$hook_write_data = 195;
	#210 spi_writer$hook_write_data = 216;
	#210 spi_writer$hook_write_data = 237;
	#210 spi_writer$hook_write_data = 2;
	#210 spi_writer$hook_write_data = 23;
	#210 spi_writer$hook_write_data = 44;
	#210 spi_writer$hook_write_data = 65;
	#210 spi_writer$hook_write_data = 86;
	#210 spi_writer$hook_write_data = 107;
	#210 spi_writer$hook_write_data = 128;
	#210 spi_writer$hook_write_data = 149;
	#210 spi_writer$hook_write_data = 170;
	#210 spi_writer$hook_write_data = 191;
	#210 spi_writer$hook_write_data = 212;
	#210 spi_writer$hook_write_data = 233;
	#210 spi_writer$hook_write_data = 254;
	#210 spi_writer$hook_write_data = 19;
	#210 spi_writer$hook_write_data = 40;
	#210 spi_writer$hook_write_data = 61;
	#210 spi_writer$hook_write_data = 82;
	#210 spi_writer$hook_write_data = 103;
	#210 spi_writer$hook_write_data = 124;
	#210 spi_writer$hook_write_data = 145;
	#210 spi_writer$hook_write_data = 166;
	#210 spi_writer$hook_write_data = 187;
	#210 spi_writer$hook_write_data = 208;
	#210 spi_writer$hook_write_data = 229;
	#210 spi_writer$hook_write_data = 250;
	#210 spi_writer$hook_write_data = 15;
	#210 spi_writer$hook_write_data = 36;
	#210 spi_writer$hook_write_data = 57;
	#210 spi_writer$hook_write_data = 78;
	#210 spi_writer$hook_write_data = 99;
	#210 spi_writer$hook_write_data = 120;
	#210 spi_writer$hook_write_data = 141;
end
 // for en_regs 

initial begin
	#1000020 $finish;
end
initial begin
	$dumpfile("tb$top.INST_counter.vcd");
	$dumpvars(0, testbench);
end
endmodule
